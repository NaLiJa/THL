���Z     @  8   I�      �   &                                       
    w                                                    !   �   �6 	   ,          � Project@Options� -�   !�     7   \+ 	   -          � File@@Version2.1  � 1.1     (                                                          1   f   TOPIC VERSION OBJARRAY BROWSE_SEQUENCE BUILD_TAG CONTEX    link viewHandles 7                                            _ISECT_iterator _AE_Sorter _AE_mark _SysInfoFlags _outside_   Metafile VbPicture VbVarArray VeRec ViewEngine WinImage _AE   r VB_Historian VB_View VbCurrency VbDibBitmap VbFixArray Vb	   ng SystemDatabase TextFileDatabase TrashCollector TreeWalke
   Real RecordMark RuleSpecifier SchemaEngine SmartString Stri   adStream NamedData NamedMonad NilMonad Number Presentation    Dictionary Integer LogStream Monad MonadArray MonadFile Mon   tion Bcd36 Boolean ClassDesc ClassMethod ComboElement Date    Set AdRec AeAccessSet AgilityDatabase ArrayDatabase Associa   ]  YAccessCombo AccessEngine AccessItem AccessRule Accessh �                   .       ,       )       8       	�     T�     W,     X�     Z�     [�     \J     ]�     ^~     _�     `I     a^     b�     cl     m�     t�     u�     v�     w                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      �0    !� BuildAll!� 0!� Inhalt!�$ � 1996 Stefan Meier, THL-Hi#   or /Link /Macro /Play /popup /Just L /Text Der THL-Editor!��   l /L /Jump Wo gibt es... /Link /Macro /Play /popup /Just L �   192,192,192), 0!�3 "Index", ( 511, 0, 511, 1023), , , (192,$   , (192,192,192), 0!�4 "Glossary", ( 0, 0, 511, 1023), , , (%    511), , , (192,192,192), 0!�. "", ( 0, 511, 1023, 511), , &   4, 64, 832, 832), , , (192,192,192), 0!�, "", ( 0, 0, 1023,'   . "The Hint Library 1.0", , , , (192,192,192), 0!�- "", ( 6(   �  �4 	   -          � F1ProjectWindowsR-�  L !�    �  !�  !�  !�  !�  !�                                      *     !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !+   �   �� 	   -          � F1ProjectButtonsZ -�   !�O  �: Bild-Anzeigefenster.,(Global), 0,<Das Bildanzeige Fenste-   7  ۬ 	   .          � F1ProjectGlossary-�   !   � 0!� 0!� No!�  !� The Hint Library 1.0!� 1!�  !�  !� /   lfe 1.0.1!�  !�  !� E:\WORK\HINT_R~1\APP.ICO!� 0!�  !�  !"    T_STRING HELP_MACRO KEYWORDS TOPIC_TITLE NOTE              A    None , !�F Title , Arial ,  18 ,  120 ,  250 ,  40 ,  40 ,2   le , Arial ,  18 ,  120 ,  250 ,  40 ,  40 ,  0 , -1 ,  0 ,3   8 ,  120 ,  250 ,  40 ,  40 ,  0 , -1 ,  0 , None , !�F Tit4    ,  40 ,  40 ,  0 , -1 ,  0 , None , !�F Title , Arial ,  15    1 , -1 ,  0 , None , !�F Title , Arial ,  18 ,  120 ,  2506    Title , Times New Roman ,  24 ,  120 ,  250 ,  40 ,  40 , 7   @'  3 	 	  ,          � F1ProjectStyle2'-�  � !�P:     � Inhaltsverzeichnis�� Q�     �  �� 	r  _-�   !;   �% /H /Just L /Text The Hint Library 1.0!�$ /T /Just L /Tex<   t  Inhaltsverzeichnis!�
 /N /Just L!� /P /Just L /Text !�T=    /L /Jump Einleitung /Link /Macro /Play /popup /Just L /Tex>   t Einleitung und �berblick!�\ /L /Jump Bedienung /Link /Mac?   ro /Play /popup /Just L /Text Allgemeine Hinweise zur Bedie@   nung!�Y /L /Jump Der THL Reader /Link /Macro /Play /popup /"   Just L /Text THL Hinweis-Dateien lesen!�J /L /Jump Der Edit�P     0 , -1 ,  0 , None , !�R Paragraph , MS Sans Serif ,  10 Q   one , !�L Sub Heading , Arial ,  12 ,  180 ,  250 ,  40 ,  B    , Arial ,  12 ,  180 ,  250 ,  40 ,  20 ,  0 , -1 , -1 , NC    ,  250 ,  60 ,  20 ,  0 , -1 ,  0 , None , !�L Sub HeadingD   20 ,  0 , -1 ,  0 , None , !�H Heading , Arial ,  12 ,  180E    , None , !�H Heading , Arial ,  12 ,  180 ,  250 ,  60 ,  F   ding , Arial ,  12 ,  180 ,  250 ,  60 ,  20 ,  0 , -1 ,  0G   2 ,  180 ,  250 ,  60 ,  20 ,  0 , -1 ,  0 , None , !�H HeaH     60 ,  20 ,  5 , -1 ,  0 , None , !�H Heading , Arial ,  1I    None , !�R Heading , Times New Roman ,  24 ,  180 ,  250 ,J   ph , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 ,K    180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�J ParagraL     60 ,  0 ,  0 ,  0 , None , !�J Paragraph , Arial ,  10 , M    , None , !�J Paragraph , Arial ,  10 ,  180 ,  250 ,  20 ,N   raph , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0O   ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�J Parag`   20 ,  0 , -1 , -1 , None , !�L Sub Heading , Arial ,  12 , a    60 ,  0 ,  0 ,  0 , None , !�N Mono Spaced , Courier ,  10R   ne , !�N Mono Spaced , Courier ,  10 ,  180 ,  250 ,  20 , S   Courier ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , NoT    250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�N Mono Spaced , U     0 ,  0 , None , !�N Mono Spaced , Courier ,  10 ,  180 , V    Jump Label , Arial ,  10 ,  180 ,  250 ,  20 ,  20 ,  10 ,W     10 ,  180 ,  250 ,  20 ,  20 ,  10 ,  0 ,  0 , None , !�LX    20 ,  20 ,  10 ,  0 ,  0 , None , !�L Jump Label , Arial ,Y   ,  0 , None , !�L Jump Label , Arial ,  10 ,  180 ,  250 , Z   p Label , Arial ,  10 ,  180 ,  250 ,  20 ,  20 ,  10 ,  0 [    ,  180 ,  250 ,  20 ,  20 ,  10 ,  0 ,  0 , None , !�L Jum\    ,  20 ,  0 , -1 , -1 , None , !�L Jump Label , Arial ,  12]    , None , !�L Sub Heading , Arial ,  12 ,  180 ,  250 ,  40^   ding , Arial ,  12 ,  180 ,  250 ,  40 ,  20 ,  0 , -1 , -1_    180 ,  250 ,  40 ,  20 ,  0 , -1 , -1 , None , !�L Sub Heap    ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�N Monoq   10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�R Bib   60 ,  0 ,  0 ,  0 , None , !�Q Bitmap Paragraph , Arial ,  c    !�Q Bitmap Paragraph , Arial ,  10 ,  180 ,  250 ,  20 ,  d   ial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None ,e    20 ,  60 ,  0 ,  0 ,  0 , None , !�Q Bitmap Paragraph , Arf    None , !�Q Bitmap Paragraph , Arial ,  10 ,  180 ,  250 , g   ph , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 ,h    250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�Q Bitmap Paragrai   ,  0 ,  0 ,  0 , None , !�H Footnote , Arial ,  8 ,  180 , j   None , !�H Footnote , Arial ,  8 ,  180 ,  250 ,  20 ,  60 k   te , Arial ,  8 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , l     180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�H Footnom   0 ,  60 ,  0 ,  0 ,  0 , None , !�H Footnote , Arial ,  8 ,n    ,  0 , None , !�H Footnote , Arial ,  8 ,  180 ,  250 ,  2o    Spaced , Courier ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0�   tmap Jump Label , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  �   �R Enumerated Bullet , Arial ,  10 ,  180 ,  250 ,  20 ,  6r   l ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !s    ,  60 ,  0 ,  0 ,  0 , None , !�R Enumerated Bullet , Ariat    ,  0 , None , !�G Bullet , Arial ,  10 ,  180 ,  250 ,  20u   �G Bullet , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0v   l ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !w     250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�G Bullet , Ariax   60 ,  0 ,  0 ,  0 , Box , !�G Bullet , Arial ,  10 ,  180 ,y   0 , None , !�F Bullet , Arial ,  10 ,  180 ,  250 ,  20 ,  z   Label , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  {   ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�R Bitmap Jump |   0 ,  0 , None , !�R Bitmap Jump Label , Arial ,  10 ,  180 }   Jump Label , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  ~    180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�R Bitmap    0 ,  0 ,  0 , None , !�R Bitmap Jump Label , Arial ,  10 , �   0 ,  0 ,  0 ,  0 , None , !�R Enumerated Bullet , Arial ,  �    ,  10 ,  440 ,  250 ,  10 ,  10 ,  0 ,  0 ,  0 , None , !��     10 ,  10 ,  0 ,  0 ,  0 , None , !�M Outline Leaf , Arial�     0 , None , !�M Outline Leaf , Arial ,  10 ,  440 ,  250 ,�   ne Leaf , Arial ,  10 ,  440 ,  250 ,  10 ,  10 ,  0 ,  0 ,�   ,  180 ,  250 ,  10 ,  10 ,  0 ,  0 ,  0 , None , !�M Outli�   0 ,  0 ,  0 ,  0 , None , !�O Outline Branch , Arial ,  10 �   , !�O Outline Branch , Arial ,  10 ,  180 ,  250 ,  10 ,  1�   rial ,  10 ,  180 ,  250 ,  10 ,  10 ,  0 ,  0 ,  0 , None �    ,  10 ,  10 ,  0 ,  0 ,  0 , None , !�O Outline Branch , A�     0 , None , !�O Outline Branch , Arial ,  10 ,  180 ,  250�    Branch , Arial ,  10 ,  180 ,  250 ,  10 ,  10 ,  0 ,  0 ,�    180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�O Outline�   0 ,  0 ,  0 , None , !�R Enumerated Bullet , Arial ,  10 , �   umerated Bullet , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  �   10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�R En�   M Outline Leaf , Arial ,  10 ,  440 ,  250 ,  10 ,  10 ,  0�   tter Label , Arial ,  12 ,  180 ,  250 ,  20 ,  60 ,  0 , -�   180 ,  250 ,  20 ,  60 ,  0 , -1 ,  0 , None , !�S Index Le�   , -1 ,  0 , None , !�S Index Letter Label , Arial ,  12 ,  �    Letter Label , Arial ,  12 ,  180 ,  250 ,  20 ,  60 ,  0 �   ,  180 ,  250 ,  20 ,  60 ,  0 , -1 ,  0 , None , !�S Index�    0 , -1 ,  0 , None , !�S Index Letter Label , Arial ,  12 �   dex Letter Label , Arial ,  12 ,  180 ,  250 ,  20 ,  60 , �   10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�S In�   50 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�E Line , Arial ,  �    ,  0 ,  0 ,  0 , None , !�E Line , Arial ,  10 ,  180 ,  2�   0 , None , !�E Line , Arial ,  10 ,  180 ,  250 ,  20 ,  60�    Line , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  �   ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�E�     250 ,  10 ,  10 ,  0 ,  0 ,  0 , None , !�E Line , Arial �    ,  0 ,  0 , None , !�M Outline Leaf , Arial ,  10 ,  440 ,��   1 ,  0 , None , !�F Index , Arial ,  10 ,  180 ,  250 ,  20�    60 ,  0 ,  0 ,  0 , None , !�I Glossary , Arial ,  10 ,  1�    , None , !�I Glossary , Arial ,  10 ,  180 ,  250 ,  20 , �   abel , Arial ,  12 ,  180 ,  250 ,  20 ,  60 ,  0 , -1 ,  0�   0 ,  20 ,  60 ,  0 , -1 ,  0 , None , !�V Glossary Letter L�   None , !�V Glossary Letter Label , Arial ,  12 ,  180 ,  25�   l , Arial ,  12 ,  180 ,  250 ,  20 ,  60 ,  0 , -1 ,  0 , �     20 ,  60 ,  0 , -1 ,  0 , None , !�V Glossary Letter Labe�   e , !�V Glossary Letter Label , Arial ,  12 ,  180 ,  250 ,�    Arial ,  12 ,  180 ,  250 ,  20 ,  60 ,  0 , -1 ,  0 , Non�   0 ,  60 ,  0 ,  0 ,  0 , None , !�V Glossary Letter Label ,�    0 ,  0 , None , !�F Index , Arial ,  10 ,  180 ,  250 ,  2�   , !�F Index , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 , �   rial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None �   80 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�F Index , A�    ,  60 ,  0 ,  0 ,  0 , None , !�F Index , Arial ,  10 ,  1�   80 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�I Glossary �   ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�D Bar ,�    ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�D Bar , Arial ,  10 �   ,  0 ,  0 ,  0 , None , !�D Bar , Arial ,  10 ,  180 ,  250�   0 , None , !�D Bar , Arial ,  10 ,  180 ,  250 ,  20 ,  60 �   D Bar , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  �    ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !��     250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�F Image , Arial�   60 ,  0 ,  0 ,  0 , None , !�F Image , Arial ,  10 ,  180 ,�    0 , None , !�F Image , Arial ,  10 ,  180 ,  250 ,  20 ,  �    Image , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 , �   ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�F�    250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�F Image , Arial �     0 ,  0 ,  0 , None , !�I Glossary , Arial ,  10 ,  180 , �   ne , !�I Glossary , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,�   , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , Noj�    Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , Non�   ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,�   1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  �   e , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !��   !�;  , Arial ,  10 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 , Non�    ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , �   0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0�    0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  �   ,  0 ,  0 ,  0 , None , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 , �    ,  0 ,  0 , None , !�;  , Arial ,  10 ,  0 ,  0 ,  0 ,  0 �   ne , !�F Table , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0�   , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , No�     180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�F Table �    20 ,  60 ,  0 ,  0 ,  0 , None , !�F Table , Arial ,  10 ,�   ,  0 ,  0 , None , !�F Table , Arial ,  10 ,  180 ,  250 , �   e , !�F Table , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 "�     0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�;  , Arial ,  10 ,�    0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 , None , !�1  ,  ,  0 ,  0�    0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�;  , Arial ,  10 , �     0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 , �     ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,�    , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1�   �;  , Arial ,  10 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 , None�   ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�    ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 �   0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0�     0 ,  0 ,  0 , None , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  �     0 ,  0 ,  0 ,  , !�;  , Arial ,  10 ,  0 ,  0 ,  0 ,  0 ,�   ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,�    ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 �   0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0�     0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 , None , !�1  ,  ,  0 ,  ��    ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 �   a normalerweise nur als Textdatei verf�gbar, der eigentlich�    oder weniger vollst�ndige Aufzeichnungen gibt, die aber, d�   spekt war, da� es an verschiedenen Stellen im Internet mehr�   r�nglich war dieses Programm nur dazu gedacht, die INVISICL�   UES(TM) zu den alten INFOCOM-Adventures in elektronischer F�   orm wiederaufzubereiten, um zu verhindern, da� diese Inform�   ationen vielleicht f�r immer verloren gehen. Ein weiterer Am  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�   Jump /Link /Macro /Play /Popup /Just L /Text !�F /L /Jump R�   /Text Wo gibt es die THL-Software und THL-Dateien ?!�1 /L /�   192,192), 0!�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  9   	  � 1000   �  ��7i     � �berblick;Inhalt;�� B�        0 ,  0 ,  0 ,  , !�                                       �     0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 , �   ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,   en Idee dieser Hinweissammlungen nicht gerecht werden. Die   puterspiele !). Um f�r m�glichst viele Menschen dieses Prog�   e zur Verf�gung zu stellen (und nicht nur unbedingt f�r Com�    aufgefordert, anderen Leuten seine besten Tips und Hinweis�   , eine Hinweis-Bibliothek aufzubauen und jeder wird hiermit�   ssammlungen anzulegen. Das nunmehr verfolgte Ziel soll sein�   ignet ist, sondern auch die M�glichkeit bietet, neue Hinwei�   ger�ckt, das nicht nur zum Lesen solcher Hinweisdateien gee�   nn immer mehr der Gedanke an ein System in den Vordergrund �   nehmen will.����Bei der Entwicklung dieses Programms ist da�   nd man selber dosieren kann, wieviel Hilfe man in Anspruch �   ich raubt, indem man in einer Komplettl�sung zuviel sieht u�   sammlungen ist, da� man sich den Spielspa� nicht versehentl�   de) Hinweise zu geben. Der gro�e Vorteil an solchen Hinweis�   blemstellen in den Textadventures (in der Pr�zision steigen�   Idee hinter den InvisiClues(tm) war es zu verschiedenen Pro�  ramm nutzbar zu machen, sollen auch m�glichst viele Sprache  cht m�glich sein. Zur Zeit begegnen Ihnen im Reader folgend  t ausw�hlen. Das versehentliche Lesen von Hinweisen soll ni  en Sie Informationen nur lesen k�nnen, wenn Sie sie explizi  e zur Verf�gung stehenden Hinweise zum Lesen an. Dabei werd  eser bietet Ihnen, normalerweise nach Themen gegliedert, di  Teilen.  Da ist zum einen der Reader, der "Lese"-Teil. Di  zum Programm selber:��Es besteht im  wesentlichen aus zwei   inen Umst�nden kommerziell genutzt werden darf.����Und nun 	  lich dem Sammeln von Informationen dienen soll und unter ke
   soll hier nochmal betont werden, da� das System ausschlie�  te, damit wir das weitere Vorgehen besprechen k�nnen.����Es  usammenzustellen. In diesem Falle kontaktieren Sie mich bit  erkl�ren w�rde, ein weiteres Sprachpaket f�r das Programm z  n. Ich w�rde mich also sehr freuen, wenn sich jemand bereit  n von der Oberfl�che und der Online-Hilfe unterst�tzt werde   e��Hinweistypen: Texte, Bilder und Multimediadateien( z.B. !  und JPEG-Dateien verwendet. Zu erreichen unter:��Meister@rz  MPICVIEW-Projekt werden von mir zur Anzeige von  PCX-,TGA-   s Meier��Alen Tomasic����Detlef Meister. Teile seines   �  	  � 2000   �  ��;�   =  �8 Sprachdateien;Sprachen;  Hinweisdateien;Infocom;�berblick;�� F�     �
 Einleitung  �� U�     �  �� 	�C  z-�   !�) /T /Just L /Text Einl�   eitung und �berblick!�
 /N /Just L!�5/P /Just L /Text Ursp  ation;Danksagung;�� B�     �
 Referenzen�� Q�     �    �� 	��  -�   !� /T /Just L /Text Referenzen!�
 /N /Ju  st L!��/P /Just L /Text Autor: Stefan Meier����Folgenden   Personen gilt mein besonderer Dank:����Beta-Tester:��Klau�  n!�P /L /Jump Lizenzvertrag /Link /Macro /Play /popup /Just  eferenzen /Link /Macro /Play /popup /Just L /Text Referenzew  esen.��Der andere Teil ist der Editor, der Ihnen die M�gl  MIDI, AVI,...)��Weiteres finden Sie unter Hinweis-Dateien-lj0  .fhtw-berlin.de����Allen Ex-Infocomlern, die mit Ihren Text#  migung entbindet den H�ndler nicht von den anderen Pflichte$  n, die sich aus diesem Vertrag ergeben.����Mein besonderer %  Dank gilt Detlef Meister f�r sein Freeware-Projekt MPICVIEW&  .��Dieses Programm nutzt Teile dieses Projektes zum Anzeige'  n von JPEG, TARGA und PCX-Dateien.��Sie erreichen Detlef Me(  ister unter;��Meister@rz.fhtw-berlin.de�� ��Kontaktadresse)  :��Stefan Meier, Erfstr. 65, D-52249 Eschweiler, Germany��*  AOL:��SMeier7777��E-Mail:��SMeier7777@aol.com��Stefan.M    eier@post.rwth-aachen.de  
� �                               �                                                            L  �L�� 
X - 4 M     � Topic@Einleitung  �      �    �    �  ��;�   1  �, Autor;Borland Delphi;Inform      
� �                                                    .  int Library 1.0 wurde mit Borland Delphi 2.0 entwickelt.��/  adventures Computergeschichte geschrieben haben.������The H""   des Programms aufh�ren.��Das Widerrufen der Vertriebsgeneh3   einer besonderen schriftlichen Genehmigung.��Kein H�ndler 4  darf mehr als 12 DM (oder den entsprechenden Betrag in ande5  ren W�hrungen, z.B. $8 US) f�r die Verbreitung dieses Progr6  amms verlangen.����Alle THL-Dateien eines H�ndlers m�ssen a7  uf eine m�glichst kleine Menge Disketten verteilt werden. D8  ie Verteilung mittels einer unnat�rlich gro�en Menge Disket9  ten ist VERBOTEN.��F�r solche Disketten, auf denen THL-Date:  ien vertrieben werden, d�rfen unter keinen Umst�nden mehr a;  ls 12 DM (oder der entsprechende Betrag in anderen W�hrunge<  n, z.B. $8 US) verlangt werden.��Diese Bedingungen gelten s=  owohl f�r die Verbreitung dieses Programms, als auch f�r al>  le THL-Dateien, die von anderen Autoren erstellt werden.���?  �Die Genehmigung zur Verteilung des Programms kann schriftl@  ich widerrufen werden. Sp�testens 30 tage nach dem Ausstell1  ungsdatum des Widerrufs, mu� der H�ndler mit der Verteilung�2  der Verbreitung �ber "Magazin-CDs" oder "Magazin-Disketten"C  , die aus der direkten oder indirekten Nutzung des ProgrammD  s entstehen, auch dann nicht, wenn der Autor auf m�gliche SE  ch�den durch die Nutzung des Programmes hingewiesen worden F  ist. ����Wenn Sie beabsichtigen, mit dem Programm THL-DateiG  en zu erstellen und zu verbreiten. sollten Sie mir mitteileH  n, welches Projekt sie vorhaben und zuerst bei mir anfragenI  , ob jemand anders gerade an einem THL-File zu dem jeweiligJ  en Thema schreibt. Obwohl das Programm unentgeldlich benutzK  t werden darf, ist es unter KEINEN UMST�NDEN ERLAUBT, f�r "L  eigene" THL-Files in irgendeiner Form Geb�hren zu verlangenM  . Wenn Sie Ihre THL-Dateien zur Verf�gung stellen wollen, sN  ollten Sie mir eine Kopie zukommen lassen. Der einfachste WO  eg ist, die Datei an der unten angegebenen FTP-Adresse abzuP  legen. �� ��Die Verbreitung �ber Warenh�user bedarf einer bA  esonderen schriftlichen Genehmigung.��Ebenso bedarf es bei �B  Stefan Meier, tr�gt in keinem Falle die Haftung f�r Sch�denS  n und m�ssen alle Kopien davon l�schen.��Dieses urheberrechT  tllich gesch�tzte Programm wird als "Freeware" vertrieben. U  Sie d�rfen das Programm unentgeldlich benutzen und an anderV  e weitergeben.��Alle Rechte an diesem Programm geh�ren StefW  an Meier und werden durch das Urheberechtsgesetz der BundesX  republik Deutschland und internationale��Abkommen gesch�tztY  . Daher mu� das Programm wie anderes gesch�tztes Material bZ  ehandelt werden (z.B. B�cher und Tontr�ger).����Dieses Prog[  ramm darf nicht vermietet werden. Au�erdem ist es nicht erl\  aubt, das Programmpaket zu ver�ndern, zu �bersetzen, zu dis]  sassemblieren oder zu decompilieren.��Wenn Sie eine der Bed^  ingungen dieses Vertrages verletzen, erlischt automatisch I_  hr Nutzungsrecht f�r dieses Programm und Sie m�ssen alle Ko`  pien l�schen.����Das Programm und die Dokumentation werden Q  so zur Verf�gung gestellt, "wie sie sind", d.h. der Autor, R  t einverstanden sind, d�rfen Sie das Programm nicht benutzec  ink E:\WORK\HINT_R~1\HELPFILE\EDITOR~1.BMP /Just L /Text Mid  t Editor - Neue Hinweisdatei erzeugen  �ffnen Sie das Edie  torfenster, um eine neue THL-Datei zu erzeugen��Mit Editorf   - Hinweisdatei editieren �ffnen Sie den Editor und sehen g  ein Dateiauswahlfenster, um eine vorhandene Datei zum Ver�nh  dern auszuw�hlen!��/R /Link E:\WORK\HINT_R~1\HELPFILE\SPRAi  CH~1.BMP /Just L /Text Mit Sprache - Sprache w�hlen �ffnej  n Sie einen Dialog, in dem Sie ein Sprachpaket ausw�hlen k�k  nnen. Standardm��ig wird mit diesem Programm das deutsche S�  prachpaket mitgeliefert. Zus�tzliche Pakete k�nnen einfach -  �  ���� 
m - 4 I     � Topic@Referenzen  �    �   !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�o  enzvertrag!�
 /N /Just L!��/P /Just L /Text Bitte lesen Sip  e diesen Lizenzvertrag komplett bevor Sie dieses Programm ba  enutzen. Wenn Sie mit den Bedingungen dieses Vertrages nich�b  der.��Mit Beenden verlassen Sie The Hint Library!�</R /Ls  en Sie unter Der THL-Editor.!�� /R /Link E:\WORK\HINT_R~1\Ht  ELPFILE\EXISTF~1.BMP /Just L /Text Hiermit �ffnen Sie den Eu  ditor, um eine bereits existierende Datei zu ver�ndern!�j /v  R /Link E:\WORK\HINT_R~1\HELPFILE\HELP.BMP /Just L /Text Miw  t diesem Knopf rufen Sie diese Hilfedatei auf.!�� /R /Link x  E:\WORK\HINT_R~1\HELPFILE\INFO.BMP /Just L /Text Hiermit �fy  fnen Sie ein Informationsfenster, in dem Sie unter anderem z  die Programmversion und Kontaktadressen finden!�^ /R /Link {  E:\WORK\HINT_R~1\HELPFILE\EXIT.BMP /Just L /Text Hiermit be|  enden Sie The Hint Library!�& /H 2 /Just L /Text Die Progra}  mm-Men�s:!� /H 2 /Just L /Text !�5/R /Link E:\WORK\HINT_R~  ~1\HELPFILE\DATEIM~1.BMP /Just L /Text Mit Datei �ffnen w  �hlen Sie eine Hinweissammlung aus und �ffnen den "Reader"��  �Mit Datei �ffnen (�ber Titel)... w�hlen Sie ein Hinweissq  ammlung nach ihrem behandelten Titel aus und �ffnen den Rea"r  ng des Editors und zum Erstellen von Hinweissammlungen find�  em Reader finden Sie unter THL-Hinweis-Dateien lesen!�� /R �  ingestellte Sprache beim n�chsten Start automatisch wieder �  Spracheinstellung speichern k�nnen Sie bestimmen, ob die e�  e mich bitte, um das weitere Vorgehen abzusprechen. ��Mit �   Verf�gung stellen k�nnten. In diesem Falle kontaktieren Si�  sehr dar�ber freuen, wenn Sie mir ein neues Sprachpaket zur�  chauen Sie bitte auf der THL-Homepage nach. Ich w�rde mich �  zu diesem Programm hinzugef�gt werden.F�r andere Sprachen s�  /Link E:\WORK\HINT_R~1\HELPFILE\VOPEN.BMP /Just L /Text Auc�  h hiermit k�nnen Sie eine THL-Datei zum Lesen �ffnen, aller�  dings sehen Sie hier nicht die Dateinamen, sondern die Tite�  l der Hinweissammlungen.!�� /R /Link E:\WORK\HINT_R~1\HELPF�  ILE\NEWFILE.BMP /Just L /Text Hiermit �ffnen Sie den Editor�     ���� 
W ) 0 I     � Topic@Inhalt  �    �  �  , um eine neue THR-Datei zu erstellen. HInweise zur Bedienu"�  ne THL-Datei zum "Hinweis-Lesen". Hinweise zum Umgang mit d�  a-�   !� /T /Just L /Text THL-Dateien!�
 /N /Just L!�/�  �     � Was sind THL Dateien...�� ^�     �  �� 	�K  �  eien;Hinweise;Bilder;Formate;THL-Dateien;THR-Dateien;�� O�  ..  �    �    �    �  ��H�   H  �C Multimedia-Dat�  tehen sie?!�| /L /Jump Eigenentwicklung von Hinweissammlung�  en /Link /Macro /Play /popup /Just L /Text Die Entwicklung �  eigener THL-Dateien.!�d /L /Jump Die Bedienung des Editors �  /Link /Macro /Play /popup /Just L /Text Die Bedienung des E�  n�s;�� E�     �	 Bedienung�� T�     �  �� 	��  �-��     !�' /T /Just L /Text Hinweise zur Bedienung!�
 /N /Just�   L!�S /P /Just L /Text Wenn Sie The Hint Library starten, s�  ehen Sie das folgende Fenster:!�3 /I /Link E:\WORK\HINT_R~1�  \HELPFILE\MAIN.BMP /Just L!� /H /Just L /Text !�( /H 2 /Ju�  st L /Text Bedeutung der Kn�pfe:!�� /R /Link E:\WORK\HINT_R�  ~1\HELPFILE\OPENBTN.BMP /Just L /Text Hiermit �ffnen Sie ei�  P /Just L /Text THL-Dateien sind Bin�rfiles, die Texte, Bil�  erschiedene Themen. Ein Thema enth�lt entweder Unterthemen �   /Just L /Text Normalerweise enth�lt eine Hinweissammlung v�  �2 /H 1 /Just L /Text Der Aufbau von THR/THL-Dateien:!�� /P�  n der Editordaten in eine THL-Datei!� /H 1 /Just L /Text !�   eine Kopie der THR-Datei !!!!�= /B /Just L /Text �bersetze�  en.��Wenn Sie eigene Dateien entwerfen, verwahren Sie immer�  G: THL-Dateien k�nnen nicht mehr im Editor bearbeitet werd�  en gespeichert, allerdings ohne sie zu �bersetzen.��ACHTUN�   SEHR EMPFOHLEN !). In einer THR-Datei werden die Editordat�  /B /Just L /Text Ggf. Abspeichern der Daten als THR-Datei (�  r Hinweise und Benennen von Bildern u.�. mit dem Editor!�D�  teien verl�uft wie folgt:!�U /B /Just L /Text Eingeben alle�   dieses Programms.��Die prinzipielle Entstehung von THL-Da�  ht mit einem Texteditor lesbar, sondern nur mit dem Reader�  der und Multimediadateien enthalten. Diese Dateien sind nic��  ODER Hinweise. Hinweise und Themen k�nnen nicht auf der gle�  Play /popup /Just L /Text Was sind THL-Dateien und wie ents�  ��Thema2 ---> Unterthema1, Hinweise1..9 ( NICHT M�GLICH )���  e Kombination ist nicht m�glich:��Thema1 ---> Hinweise 1..3�  ema1,Unterthema2��Thema3 ---> Bild, Hinweis 1..6����Folgend�  st m�glich:��Thema1 ---> Hinweise 1..3��Thema2 ---> Unterth�  �'/P /Just L /Text Zwei Beispiele:��Folgende Kombination i�  sicher, da� jeder diese Hinweise lesen/ansehen/h�ren kann.!�  eitere Formate unterst�tzt, allerdings ist dann nicht mehr �  t�tzt werden WAV, AVI, MIDI, MOV. Prinzipiell werden auch w�  en versehen.!�� /B /Just L /Text Multimedia-Dateien, unters�  e aus Bildern definieren und diese mit eigenen Beschreibung�   Targa��Besonderheiten: Sie k�nnen mit dem Editor Auschnitt�  st L /Text Bilder, unterst�tzte Formate: Bitmap, JPeg, PCX,�  / /B /Just L /Text Texte ( ein- oder mehrzeilig )!�� /B /Ju�  ichen Ebene liegen. Folgende Typen von Hinweisen gibt es:!��   /Just L!�t /L /Jump Was sind THL Dateien... /Link /Macro /�  klaren, fragen Sie beim Inhaber der Urheberrechte um Erlaub�  nis.!�1/B /Just L /Text Verbreiten sollten Sie normalerwei�  se nur die THL-Datei, damit au�er Ihnen keine die Daten ver�  �ndern kann. WICHTIG: Behalten Sie aber immer eine Kopie �  der THR-Datei, da sie sonst auch selber Ihre Daten nicht me�  hr �ndern k�nnen. EINE THL-DATEI KANN NICHT MEHR IM EDITOR �  VER�NDERT WERDEN !!�E/B /Just L /Text Lassen Sie mir eine �  Kopie Ihrer THL-Datei zukommen. Am einfachsten geht dies, i�  p://members.aol.com/thlhome/incoming��Sie k�nnen mir auch �  eine Diskette per Post schicken, oder mir eine Adresse im I+  nternet benennen, unter der die Datei erh�ltlich ist  
� �  ndem Sie die Datei an die folgende ftp-Adresse senden:��ft    ditors  
� �                                             �  ateien,editieren;�� F�     �
 Der Editor�� U�     �  �  �� 	�P  �-�   !� /T /Just L /Text Der THL-Editor!�
 /Nj�  Form zu �bertragen. Sind Sie sich �ber die Rechtslage im un�   sollten Sie folgende Hinweise beherzigen:!�d/B /Just L /T�  ext Bevor Sie mit Ihrer Arbeit beginnen, kontaktieren Sie m�  ich, um zu erfragen, ob schon jemand anderes an einer Datei�   zu Ihrem Spiel / Thema arbeitet. Dies soll einerseits verh�  indern, da� Arbeit unn�tigerweise doppelt gemacht wird und �  andererseits gibt es mir die M�glichkeit, einen �berblick ��  ber die Entwicklung des THL-Projekts zu bewahren!�� /B /Jus�  t L /Text �berlegen Sie sich eine Gliederung f�r Ihre Hinwe�  issammlung. Wo treten Fragen auf ? Wo kann man Sinnabschnit�  te abgrenzen? Wo ist Bildmaterial hilfreich ?!�� /B /Just L�   /Text Vergleichen Sie Ihre L�sungswege, wenn m�glich, mit �  anderen L�sungen, um Fehler oder Auslassungen zu vermeiden.�  !�'/B /Just L /Text Bitte achten Sie darauf, da� Sie keine�   Urheberrechte verletzen. So ist es normalerweise nicht erl�  aubt, kommerziell vertriebene "Hintbooks" in elektronische ��  n, eigene Hinweissammlungen zu entwerfen und zu verbreiten,    :��http://members.aol.com/thlhome/index.htm  
� �        �   zus�tzliche Sprachpackete und THL-Dateien finden Sie unter�  ?!�
 /N /Just L!�� /B /Just L /Text Neue Programmversionen,�    �  �� 	��  � -�   !�  /T /Just L /Text Wo gibt es... �  teien;Neue Versionen;�� I�     � Wo gibt es ?�� X�   �    �  	  � 8000   �  ��>�   .  �) Sprachdateien;THL-Da`    !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�   L /Text Lizenzbedingungen!�; /P /Just L /Text ������The Hi�    �  	  � 7000   �  ��>�   8  �3 Benutzung, Bedingung�  en;Vertriebsbedingungen;Lizenz;�� I�     � Lizenzvertran  g�� X�     �  �� 	��  
-�   !� /T /Just L /Text Liz�   Entwicklung;Eigene Dateien;THL-Dateien;�� ^�   +  �& Eig�  enentwicklung von Hinweissammlungen�� m�     �  �� 	��    -�  	 !�0 /T /Just L /Text Entwicklung eigener THL-Date�  ien!�
 /N /Just L!�� /P /Just L /Text Wenn Sie beabsichtige#�    �  	  � 8000   �  ��>�   .  �) Sprachdateien;THL-Da  E:\WORK\HINT_R~1\HELPFILE\EDITOR.BMP /Macro /Play /Popup /J�   Bedienung des THL-Editors!�
 /N /Just L!�O /I /Jump /Link �  s�� d5    �  �� 	�  �-�   !�. /T /Just L /Text Die�  , Bedienung;Editor;�� U%    � Die Bedienung des Editor�  rmate;Dateien bearbeiten;THL-Dateien;THR-Dateien;THL-Editor�  T  P�� 
T : A V   "  � Topic@Was sind THL Dateien.�  Hinweissammlungen  �    �    �    �  ��W�   ,  �'�  rt;Autor;Titel;Themen;Bilder;Multimedia-Dateien;Hinweise;Fo�  tors  �    �  	  � 6000   �  ��J�   �  �� Schrifta�  �  4n�� 
Z < C \   $  � Topic@Die Bedienung des EdiQ  geladen wird.!��/R /Link E:\WORK\HINT_R~1\HELPFILE\HILFEM~�  �  �N�� 
w , 3 L     � Topic@Bedienung  �    ��    	  � 3000   �  ��:w   !  � Sprachen;Hauptfenster;Me    nt Library � 1996 Stefan Meier  
� �                          !�                                                        "  ust L!�P /P /Just L /Text BITTE BEACHTEN SIE DIE HINWEISE Z  �nnen Sie einen neuen Hinweis in Ihr Projekt einf�gen. Dazu  ierfenster ge�ffnet.!�� /E /Just L /Text Mit diesem Knopf k  jekt ein neues Thema hinzuf�gen. Dabei wird das Themen-Edit  ust L /Text Bei Dr�cken dieses Knopfes k�nnen Sie Ihrem Pro  m, wa Sie f�r diesen Eintrag noch einf�gen k�nnen.!�� /E /J  Element selektieren ver�ndern sich die Kn�pfe 2-5 je nachde  er jeweis selektierte Eintrag als "Besitzer". Wenn Sie ein   mediadateien. Wenn Sie neue Eintr�ge hinzuf�gen, fungiert d	  alten ENTWEDER Unterthemen ODER Hinweise,��Bilder und Multi
  pt>>>) kann nur Themen enthalten. Die einzelnen Themen enth  ersten Buchstaben des Titels. Das Hauptverzeichnis (<<<Scri  ort PIC und Multimediadateien MM. Bei Themen sehen Sie sie   ihrem Eintrag das Schl�sselwort HINT, Bilder das Schl�sselw  en Sie Ihr Projekt als Baumansicht, Hinweise enthalten vor   UM ERSTELLEN VON THL-DATEIEN !!�^/E /Just L /Text Hier seh    wird das Hinweis-Editierfenster ge�ffnet!�� /E /Just L /Te!  dern, d.h. Sie k�nnen nicht aus einem Thema einen Hinweis m  ffnet. Es ist nicht m�glich den Typ eines Eintrags zu ver�n  dern. Je nach Typ wird das entsprechende Editierfenster ge�   Mit diesem Knopf k�nnen Sie den selektierten Eintrag ver�n   manche Benutzer nicht mehr lesbar sind!�/E /Just L /Text   daran denken, da� ausgefallene Multimedia-Formate u.U. f�r  ine von den F�higkeiten Ihres Systems abh�ngen, sollten Sie  HL-Datei anw�chst. Obwohl die Multimedia-Unterst�tzung alle  n in der Regel relativ gro� sind und dementsprechend Ihre T  ge�ffnet. Bitte beachten sie hierbei, da� z.B. Video-Dateie  jekt hinzuzuf�gen. Dazu wird das Multimedia-Editierfenster    Nummer 5 erlaubt es Ihnen, Multimedia-Dateien zu Ihrem Pro   Bildbereiche definieren k�nnen..!��/E /Just L /Text Knopf  en neuen Bildeintrag zu Ihrem Projekt hinzuf�gen k�nnen und  xt Hier �ffnen Sie das Bild-Editierfenster, mit dem Sie ein�0  achen usw.!�� /E /Just L /Text Hiermit k�nnen Sie den momen1  alle Schriftarten zur Verf�gung haben, die auf Ihrem System"  stellen. Bitte beachten Sie, da� andere Benutzer evt.nicht #  rt w�hlen, die im Reader benutzt wird, um Ihren Titel darzu$  Just L /Text Mit dem Schrift-Knopf k�nnen Sie eine Schrifta%  �llt sein, damit Ihr Projekt �bersetzt werden kann.!�u/E /&  tel, der sp�ter im Reader erscheint. Dieses Feld mu� ausgef'  f�r Ihr Projekt an. Dies ist kein Dateiname, sondern der Ti(  en"!�� /E /Just L /Text In diesem Feld geben Sie den Titel )  �; /E /Just L /Text Analog zu Knopf 8 "Verschieben nach unt*  h wird werden evt. vorhandene Untereintr�ge mit verschoben!+  intrag innerhalb seiner Ebene nach oben zu verschieben. Auc,  ust L /Text Dieser Knopf gibt Ihnen die M�glichkeit einen E-  en Sie also bitte vorsichtig mit dieser Funktion !!�� /E /J.  einem Eintrag auch alle evt. vorhandenen Untereintr�ge. Sei/  tan selektierten Eintrag l�schen. ACHTUNG: Sie l�schen mit �@   installiert sind. Um unerw�nschte Effekte zu vermeiden, so3   ein. Schlie�en Sie das Fenster mit OK, wird das Thema zu I    hrem Projekt hinzugef�gt.  
� �                          �  �  	  � 5000   �  ��;�   -  �( THL-Editor;Editor;THL-Dz  ROJEKT IN JEDEM STADIUM DER ENTWICKLUNG EINE THR-DATEI ZU E5   ver�ndern wollen. ES WIRD UNBEDINGT EMPFOHLEN, VON IHREM P6  mat. Sie ben�tigen diese Datei, wenn Sie Ihr Projekt sp�ter7  n Sie einen Dialog zum Speichern Ihres Projektes im THR-For8  ojekt einzugeben!�/E /Just L /Text Mit diesem Knopf �ffne9  hnen die M�glichkeit, zus�tzliche Informationen zu Ihrem Pr:   1996 Harry Hummel.!�n /E /Just L /Text Dieses Feld gibt I;   Beispiel: Written 1996 by Harry Hummel oder Copyright �<  � ausgef�llt sein, damit das Projekt �bersetzt werden kann.=  e Informationen �ber sich als Autor an. Auch dieses Feld mu>  liefert werden.!�� /E /Just L /Text In diesem Feld geben Si?  llten Sie nur Schriftarten verwenden, die beim System mitge2   /Just L /Text Unter Text tragen Sie den Titel Ihres Themas�  weis ein. Wenn Sie das Fenster mit OK schlie�en, wird der HB  /Just L!�� /P /Just L /Text Unter Text tragen Sie Ihren HinC  E:\WORK\HINT_R~1\HELPFILE\HINTEDIT.BMP /Macro /Play /Popup D  Das Hinweis-Editierfenster!�
 /N /Just L!�Q /I /Jump /Link E  ster�� e�     �  �� 	�  9-�   !�+ /T /Just L /Text F  eingabe;Text;Hinweis;�� V�     � Das Hinweis EditierfenG  nster  �    �  	  � 5020   �  ��K�   !  � HinweisH    ?O�� 
a = D ]   %  �  Topic@Das Hinweis EditierfeK  �  ���� 
] < C \   $  � Topic@Das Themen EditierfenL  ster  �    �  	  � 5030   �  ��J~     � ThemeneiM  ngabe;Text;�� U�     � Das Themen Editierfenster�� d�N       �  �� 	��  +-�   !�* /T /Just L /Text Das Themen-P  Editierfenster!�
 /N /Just L!�P /I /Jump /Link E:\WORK\HINT_  r>!�1 Bild-Editierfenster,Das Bilder Editierfenster, 0,!�' A  _R~1\HELPFILE\TOPEDIT.BMP /Macro /Play /Popup /Just L!�� /P�  1.BMP /Just L /Text Mit Hilfe - Inhalt rufen Sie diese Hia   Sie die linke Maustaste loslassen, wird der Auschnitt IhreR  arkieren den Bildauschnitt, den Sie benennen wollen. SobaldS  aste in das Bild, halten die linke Maustaste gedr�ckt und mT  ldhinweise eintragen. Dazu klicken Sie mit der linken MaustU  seditor k�nnen Sie separate Bildausschnitte als einzelne BiV  d die jeweils behandelte Bilddatei eingetragen.  Im BereichW  ro /Play /Popup /Just L!��/P /Just L /Text Unter Datei wirX  P /I /Jump /Link E:\WORK\HINT_R~1\HELPFILE\PICEDIT.BMP /MacY   /T /Just L /Text Das Bilder-Editierfenster!�
 /N /Just L!�Z   Bilder Editierfenster�� d�     �  �� 	�%  F-�   !�*[  ten;Bilder;Fortschrittsanzeige;Bereiche;�� U�     � Das\  ster  �    �  	  � 5010   �  ��J�   5  �0 Koordina]  .  N��� 
b < C \   $  � Topic@Das Bilder Editierfenh  Der THL-Editor,(Global), 0,<Der Editor>!�' Der-THL-Editor,(    �  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�      p  r Bereichsliste hinzugef�gt. Sie m�ssen dann noch eine Bescc   /Just L /Text Das Multimedia-Editierfenster!�
 /N /Just L!d  �O /I /Jump /Link E:\WORK\HINT_R~1\HELPFILE\MMEDIT.BMP /Mace  ro /Play /Popup /Just L!�� /P /Just L /Text Unter Datei traf  gen Sie die behandelte Multimedia-Datei ein. Unter Beschreig  bung geben Sie der Datei einen Titel. Wenn Sie das Fenster �  mit OK schlie�en, wird dieser Multimedia-Eintrag zum aktuel}  Global), 0,<Der Editor>!�Q Eigene THL-Dateien erstellen,(Gl�  d sp�ter im Reader jeder eingetragene Bereich als ein einzei  ohl Sie im Editor nur einen Eintrag f�r ein Bild sehen, wirj  zu dem aktuell selektierten Thema hinzugef�gt. Beachte: Obwk  enn Sie das Fenster mit OK schlie�en, wird der Bildeintrag l  diesen eintrag nicht w�nschen, ihn aus der Liste l�schen. Wm  Sie sollten die Beschreibung hierzu �ndern, oder falls Sie n  rd automatisch das komplette Bild als Bereich eingetragen. o  hreibung hinzuf�gen. Wenn Sie eine neue Datei ausw�hlen, wi"b  edia Editierfenster�� h�     �  �� 	�`  �-�   !�. /T�  -THL-Editor. ( Bitte unbedingt lesen ! )��Nicht zu sehen isr  itor und zum Erstellen von THL-Dateien finden Sie unter Ders  PEG, TARGA, PCX) in Ihre Dateien aufnehmen.��N�heres zum Edt  Sie Multimediadateien ( Sound, Videos ) und Bilder ( BMP, Ju  komfortabel in einem Fenster erledigt. Neben Texten k�nnen v  ichkeit gibt, neue Hinweis- Dateien anzulegen. Dieses wird �  >!�5 Hinweis-Editierfenster,Das Hinweis Editierfenster, 0,!x  nweis Fenster>!�* Hinweis-Dateien-lesen,(Global), 0,<(None)�  RSTELLEN !!�k /E /Just L /Text Mit diesem Knpof �ffnen Sie y  issammlungen>!�8 Hinweis-Anzeigefenster,(Global), 0,<Das Hi{  LEN VON THL-DATEIEN,(Global), 0,<Eigenentwicklung von Hinwe|  obal), 0,<Eigenentwicklung von Hinweissammlungen>!�N ERSTEL  i  ��� 
_ @ G `   (  �# Topic@Das Multimedia Editie�  rfenster  �    �  	  � 5040   �  ��N�   *  �% Multq  imedia-Dateien;Dateibeschreibung;�� Y�   "  � Das Multim��  t der "�bersetzer", der aus Ihren "Rohdaten" eine THL-Datei�  n, �ffnet sich das Hinweis-Anzeigefenster. Anmerkung:��Da d�  inweise. Wenn Sie durch Doppelklicken einen Hinweis anw�hle�  k E:\WORK\HINT_R~1\HELPFILE\HINTPIC.BMP /Just L /Text F�r H�  der Hinweise. Diese sehen in etwa wie folgt aus:!�i/R /Lin�  ine Ebene tiefer. Dort finden Sie entweder weitere Themen o�  h�lt. Durch doppeltes Anklicken eines Themas gelangen Sie e�  n der mitte sehen Sie die Hauptthemen, welche die datei ent�  pup /Just L!�/P /Just L /Text In dem Aufz�hlungsfenster i�  /Link E:\WORK\HINT_R~1\HELPFILE\READER.BMP /Macro /Play /Po�  n einer THL-Datei sehen Sie folgendes Fenster:!�O /I /Jump �  N /Just L!�\ /P /Just L /Text Nach der �ffnen und �bersetze�   �� 	��  �-�   !� /T /Just L /Text Der THL-Reader!�
 /�  Reader;Reader;�� J�     � Der THL Reader�� Y�     � �    �  	  � 4000   �  ��?�   &  �! Hinweise lesen;THL-�  �  Z��� 
[ 1 8 Q     � Topic@Der THL Reader  �  ��  ie Hinweise einer Auswahl in der Pr�zision ansteigen, wird �  r ge�ffnet, mit dem Sie die Multimedia-datei abspielen k�nn�  en. Mit OK schlie�en Sie das Fenster. Dabei noch laufende A�  �; Multimedia-Editierfenster,Das Multimedia Editierfenster,�  ^�     �  �� 	�8  s-�   !�$ /T /Just L /Text Das Hinw�  weis;Hinweis zeigen;�� O�     � Das Hinweis Fenster�� �    �    �  	  � 4020   �  ��D�   '  �" Verdeckter Hin�  A  ���� 
` 6 = V     � Topic@Das Hinweis Fenster�  en ein Bild anw�hlen, �ffnet sich das Bild-Anzeigefenster.�  IC.BMP /Just L /Text F�r Bilder. Wenn Sie durch Doppelklick�  Kontrollfenster.!�� /R /Link E:\WORK\HINT_R~1\HELPFILE\PICP�  ine Multimedia-Datei ausw�hlen, �ffnet sich das Multimedia-�  ext F�r Multimedia-Hinweise. Wenn Sie durch Doppelklicken e�  !�� /R /Link E:\WORK\HINT_R~1\HELPFILE\MMPIC.BMP /Just L /T�  lesen wollen, bevor Sie die Hinweise 1 und 2 gelesen haben.�  eine Warnung erscheinen, wenn Sie beispielsweise Hinweis 3 ��  r Auswahl einer Multimedia-Datei wird dieses Kontrollfenste�  "Schlie�en" das Fenster zumachen. Dabei wird dieser Hinweis�  den Knopf "Hinweis zeigen" dr�cken. Danach k�nnen Sie mit  �   Sie das folgende Fenster. Um den Text zu lesen, m��en Sie �  Just L /Text Wenn Sie einen Hinweis ausgew�hlt haben, sehen�  1\HELPFILE\HINTVIEW.BMP /Macro /Play /Popup /Just L!��/P /�  eis-Fenster!�
 /N /Just L!�Q /I /Jump /Link E:\WORK\HINT_R~�  ia Fenster>!�3 Themen-Editierfenster,Das Themen Editierfens�   0,!�? Multimedia-Kontrollfenster,(Global), 0,<Das Multimed�  ~  ���� 
^ 9 @ Y   !  � Topic@Das Multimedia Fenste�  r  �    �  	  � 4030   �  ��G�   G  �B Multimedia-�  Kontrolle;Multimediadateien abspielen;Multimediaplayer;�� �  R�     � Das Multimedia Fenster�� a�     �  �� 	�u �   �-�   !�' /T /Just L /Text Das Multimedia-Fenster!�
 /N �  /Just L!�O /I /Jump /Link E:\WORK\HINT_R~1\HELPFILE\MMVIEW.�  BMP /Macro /Play /Popup /Just L!�� /P /Just L /Text Nach de�   innerhalb der momentan g�ltigen Auswahlliste als Gelesen m    inweis zum aktuell selektierten Thema hinzugef�gt.  
� �     lner Hinweis behandelt.  
� �                            �  �  �a�� 
c : A Z   "  � Topic@Das Bildanzeige Fenst�  er  �    �  	  � 4010   �  ��H�      � Fortschrit�  tsanzeige;Bilder;�� S�     � Das Bildanzeige Fenster���   b�     �  �� 	��  %-�   !�( /T /Just L /Text Das Bil�  danzeige-Fenster!�
 /N /Just L!�P /I /Jump /Link E:\WORK\HI�  ter, 0,!�- THL-Homepage nach,(Global), 0,<Wo gibt es...>!� �  NT_R~1\HELPFILE\PICVIEW.BMP /Macro /Play /Popup /Just L!�� �  /P /Just L /Text Die Anzeige unten rechts gibt den Fortschr�  itt beim Laden des Bildes an. Mit Schlie�en verlassen Sie d    as Bildanzeige-Fenster.  
� �                            �  nnen Sie das Fenster mit dem Close-Icon oben rechts schlie��  cht ist Ihnen ja inzwischen eine neue Idee gekommen), so k��  arkiert. Wollen Sie einen Hinweis doch nicht lesen (viellei    en  
� �                                                 �  um Umgang mit dem Windows Hilfesystem��Info zeigt Ihnen e�  lw�rtern suchen��Hilfe-benutzen zeigt Ihnen Erkl�rungen z�  - Suchen k�nnen Sie in der ganzen Hilfedatei nach Schl�sse�  lfedatei auf und starten im Inhaltsverzeichnis��Mit Hilfe �  �  � �� 
t 0 7 P     � Topic@Wo gibt es...  �      ...  
� �                                                �  �  ��� 
u 0 7 P     � Topic@Lizenzvertrag  �  �    ���� 
v I P e   1  �, Topic@Eigenentwicklung von     tte speichern Sie Ihr Projekt vor dem Schlie�en ! 
.> �  ei.!�e /E /Just L /Text Hiemit schlie�en Sie den Editor. Bi�  einen Dialog zum �bersetzen Ihres Projektes in eine THL-Dat      
� �                                                    4  Y  ��� 
\ - 4 M     � Topic@Der Editor  �        bspielvorg�nge werden automatisch gestoppt.  
� �            len Thema hinzugef�gt.  
� �                             �  in Fenster, dem Sie die aktuelle Programmversion, Kontaktad                                                               �                                                             �  �  ���� 
S 0 7 P     � Topic@Wo gibt es...  �                                                                     
� �                                                      �  index.htm����Viel Vergn�gen mit THE HINT LIBRARY !������  �  bers.aol.com/thlhome��oder��http://members.aol.com/thlhome/�  ost.rwth-aachen.de����The Hint Library Homepage:��ftp://mem�  l:   SMeier7777@aol.com oder��               Stefan.Meier@p�  , Erfstr. 65, 52249 Eschweiler��AOL:      SMeier7777��e-Mai�  rn o.�. erreichen Sie mich unter:��Post:       Stefan Meier�  ene THL-Dateien erstellen.����Bei Fragen, Anregungen, Fehle�   generiert.��Informationen hierzu finden Sie im Kapitel Eig�  �  �� 
d , 3 L     � Topic@Bedienung  �    �    ressen und weitere Informationen entnehmen k�nnen  
� �  