���Z     @  G   I�      /   &                                       
    �                                                    !   �   R� 	   ,          � Project@Options� -�   !�     7   \+ 	   -          � File@@Version2.1  � 1.1     (                                                          1   f   TOPIC VERSION OBJARRAY BROWSE_SEQUENCE BUILD_TAG CONTEX    link viewHandles 7                                            _ISECT_iterator _AE_Sorter _AE_mark _SysInfoFlags _outside_   Metafile VbPicture VbVarArray VeRec ViewEngine WinImage _AE   r VB_Historian VB_View VbCurrency VbDibBitmap VbFixArray Vb	   ng SystemDatabase TextFileDatabase TrashCollector TreeWalke
   Real RecordMark RuleSpecifier SchemaEngine SmartString Stri   adStream NamedData NamedMonad NilMonad Number Presentation    Dictionary Integer LogStream Monad MonadArray MonadFile Mon   tion Bcd36 Boolean ClassDesc ClassMethod ComboElement Date    Set AdRec AeAccessSet AgilityDatabase ArrayDatabase Associa   ]  YAccessCombo AccessEngine AccessItem AccessRule Accessh                   .       ,       )       8       	�     v�     {�     �     �~     �J     ��     ��     �     ��     �-     ��     ��     ��     ��     ��     ��     ��     ��     �     �     �0     �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �0    !� BuildAll!� 0!� Inhalt!�' � 1996-97 Stefan Meier, THL#   /Text Wo gibt es die THL-Software und THL-Dateien ?!�1 /L /�   Jump /Link /Macro /Play /Popup /Just L /Text !�\ /L /Jump W�   192,192,192), 0!�3 "Index", ( 511, 0, 511, 1023), , , (192,$   , (192,192,192), 0!�4 "Glossary", ( 0, 0, 511, 1023), , , (%    511), , , (192,192,192), 0!�. "", ( 0, 511, 1023, 511), , &   4, 64, 832, 832), , , (192,192,192), 0!�, "", ( 0, 0, 1023,'   . "The Hint Library 1.1", , , , (192,192,192), 0!�- "", ( 6(   �  �� 	   -          � F1ProjectWindows�-�  ] !�    �  !�  !�  !�  !�  !�                                      *     !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !+   �   �� 	   -          � F1ProjectButtonsZ -�   !�O  �: Bild-Anzeigefenster.,(Global), 0,<Das Bildanzeige Fenste-   �  `� 	   .          � F1ProjectGlossary{-�   !    !�  !� 0!� 0!� No!�  !� The Hint Library 1.1!� 1!�  !/   -Hilfe 1.1.1!�  !�  !� E:\WORK\HINT_R~1.11\APP.ICO!� 0!� "    T_STRING HELP_MACRO KEYWORDS TOPIC_TITLE NOTE              A    None , !�F Title , Arial ,  18 ,  120 ,  250 ,  40 ,  40 ,2   le , Arial ,  18 ,  120 ,  250 ,  40 ,  40 ,  0 , -1 ,  0 ,3   8 ,  120 ,  250 ,  40 ,  40 ,  0 , -1 ,  0 , None , !�F Tit4    ,  40 ,  40 ,  0 , -1 ,  0 , None , !�F Title , Arial ,  15    1 , -1 ,  0 , None , !�F Title , Arial ,  18 ,  120 ,  2506    Title , Times New Roman ,  24 ,  120 ,  250 ,  40 ,  40 , 7   @'  3 	 	  ,          � F1ProjectStyle2'-�  � !�P:   t  Inhaltsverzeichnis!�
 /N /Just L!� /P /Just L /Text !�T;    /L /Jump Einleitung /Link /Macro /Play /popup /Just L /Tex<   t Einleitung und �berblick!�\ /L /Jump Bedienung /Link /Mac=   ro /Play /popup /Just L /Text Allgemeine Hinweise zur Bedie>   nung!�Y /L /Jump Der THL Reader /Link /Macro /Play /popup /?   Just L /Text THL Hinweis-Dateien lesen!�J /L /Jump Der Edit@   or /Link /Macro /Play /popup /Just L /Text Der THL-Editor!�"   l /L /Jump Wo gibt es... /Link /Macro /Play /popup /Just L �P     0 , -1 ,  0 , None , !�R Paragraph , MS Sans Serif ,  10 Q   one , !�L Sub Heading , Arial ,  12 ,  180 ,  250 ,  40 ,  B    , Arial ,  12 ,  180 ,  250 ,  40 ,  20 ,  0 , -1 , -1 , NC    ,  250 ,  60 ,  20 ,  0 , -1 ,  0 , None , !�L Sub HeadingD   20 ,  0 , -1 ,  0 , None , !�H Heading , Arial ,  12 ,  180E    , None , !�H Heading , Arial ,  12 ,  180 ,  250 ,  60 ,  F   ding , Arial ,  12 ,  180 ,  250 ,  60 ,  20 ,  0 , -1 ,  0G   2 ,  180 ,  250 ,  60 ,  20 ,  0 , -1 ,  0 , None , !�H HeaH     60 ,  20 ,  5 , -1 ,  0 , None , !�H Heading , Arial ,  1I    None , !�R Heading , Times New Roman ,  24 ,  180 ,  250 ,J   ph , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 ,K    180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�J ParagraL     60 ,  0 ,  0 ,  0 , None , !�J Paragraph , Arial ,  10 , M    , None , !�J Paragraph , Arial ,  10 ,  180 ,  250 ,  20 ,N   raph , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0O   ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�J Parag`   20 ,  0 , -1 , -1 , None , !�L Sub Heading , Arial ,  12 , a    60 ,  0 ,  0 ,  0 , None , !�N Mono Spaced , Courier ,  10R   ne , !�N Mono Spaced , Courier ,  10 ,  180 ,  250 ,  20 , S   Courier ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , NoT    250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�N Mono Spaced , U     0 ,  0 , None , !�N Mono Spaced , Courier ,  10 ,  180 , V    Jump Label , Arial ,  10 ,  180 ,  250 ,  20 ,  20 ,  10 ,W     10 ,  180 ,  250 ,  20 ,  20 ,  10 ,  0 ,  0 , None , !�LX    20 ,  20 ,  10 ,  0 ,  0 , None , !�L Jump Label , Arial ,Y   ,  0 , None , !�L Jump Label , Arial ,  10 ,  180 ,  250 , Z   p Label , Arial ,  10 ,  180 ,  250 ,  20 ,  20 ,  10 ,  0 [    ,  180 ,  250 ,  20 ,  20 ,  10 ,  0 ,  0 , None , !�L Jum\    ,  20 ,  0 , -1 , -1 , None , !�L Jump Label , Arial ,  12]    , None , !�L Sub Heading , Arial ,  12 ,  180 ,  250 ,  40^   ding , Arial ,  12 ,  180 ,  250 ,  40 ,  20 ,  0 , -1 , -1_    180 ,  250 ,  40 ,  20 ,  0 , -1 , -1 , None , !�L Sub Heap    ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�N Monoq   10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�R Bib   60 ,  0 ,  0 ,  0 , None , !�Q Bitmap Paragraph , Arial ,  c    !�Q Bitmap Paragraph , Arial ,  10 ,  180 ,  250 ,  20 ,  d   ial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None ,e    20 ,  60 ,  0 ,  0 ,  0 , None , !�Q Bitmap Paragraph , Arf    None , !�Q Bitmap Paragraph , Arial ,  10 ,  180 ,  250 , g   ph , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 ,h    250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�Q Bitmap Paragrai   ,  0 ,  0 ,  0 , None , !�H Footnote , Arial ,  8 ,  180 , j   None , !�H Footnote , Arial ,  8 ,  180 ,  250 ,  20 ,  60 k   te , Arial ,  8 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , l     180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�H Footnom   0 ,  60 ,  0 ,  0 ,  0 , None , !�H Footnote , Arial ,  8 ,n    ,  0 , None , !�H Footnote , Arial ,  8 ,  180 ,  250 ,  2o    Spaced , Courier ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0�   tmap Jump Label , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  �   �R Enumerated Bullet , Arial ,  10 ,  180 ,  250 ,  20 ,  6r   l ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !s    ,  60 ,  0 ,  0 ,  0 , None , !�R Enumerated Bullet , Ariat    ,  0 , None , !�G Bullet , Arial ,  10 ,  180 ,  250 ,  20u   �G Bullet , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0v   l ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !w     250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�G Bullet , Ariax   60 ,  0 ,  0 ,  0 , Box , !�G Bullet , Arial ,  10 ,  180 ,y   0 , None , !�F Bullet , Arial ,  10 ,  180 ,  250 ,  20 ,  z   Label , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  {   ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�R Bitmap Jump |   0 ,  0 , None , !�R Bitmap Jump Label , Arial ,  10 ,  180 }   Jump Label , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  ~    180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�R Bitmap    0 ,  0 ,  0 , None , !�R Bitmap Jump Label , Arial ,  10 , �   0 ,  0 ,  0 ,  0 , None , !�R Enumerated Bullet , Arial ,  �    ,  10 ,  440 ,  250 ,  10 ,  10 ,  0 ,  0 ,  0 , None , !��     10 ,  10 ,  0 ,  0 ,  0 , None , !�M Outline Leaf , Arial�     0 , None , !�M Outline Leaf , Arial ,  10 ,  440 ,  250 ,�   ne Leaf , Arial ,  10 ,  440 ,  250 ,  10 ,  10 ,  0 ,  0 ,�   ,  180 ,  250 ,  10 ,  10 ,  0 ,  0 ,  0 , None , !�M Outli�   0 ,  0 ,  0 ,  0 , None , !�O Outline Branch , Arial ,  10 �   , !�O Outline Branch , Arial ,  10 ,  180 ,  250 ,  10 ,  1�   rial ,  10 ,  180 ,  250 ,  10 ,  10 ,  0 ,  0 ,  0 , None �    ,  10 ,  10 ,  0 ,  0 ,  0 , None , !�O Outline Branch , A�     0 , None , !�O Outline Branch , Arial ,  10 ,  180 ,  250�    Branch , Arial ,  10 ,  180 ,  250 ,  10 ,  10 ,  0 ,  0 ,�    180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�O Outline�   0 ,  0 ,  0 , None , !�R Enumerated Bullet , Arial ,  10 , �   umerated Bullet , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  �   10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�R En�   M Outline Leaf , Arial ,  10 ,  440 ,  250 ,  10 ,  10 ,  0�   tter Label , Arial ,  12 ,  180 ,  250 ,  20 ,  60 ,  0 , -�   180 ,  250 ,  20 ,  60 ,  0 , -1 ,  0 , None , !�S Index Le�   , -1 ,  0 , None , !�S Index Letter Label , Arial ,  12 ,  �    Letter Label , Arial ,  12 ,  180 ,  250 ,  20 ,  60 ,  0 �   ,  180 ,  250 ,  20 ,  60 ,  0 , -1 ,  0 , None , !�S Index�    0 , -1 ,  0 , None , !�S Index Letter Label , Arial ,  12 �   dex Letter Label , Arial ,  12 ,  180 ,  250 ,  20 ,  60 , �   10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�S In�   50 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�E Line , Arial ,  �    ,  0 ,  0 ,  0 , None , !�E Line , Arial ,  10 ,  180 ,  2�   0 , None , !�E Line , Arial ,  10 ,  180 ,  250 ,  20 ,  60�    Line , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  �   ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�E�     250 ,  10 ,  10 ,  0 ,  0 ,  0 , None , !�E Line , Arial �    ,  0 ,  0 , None , !�M Outline Leaf , Arial ,  10 ,  440 ,��   1 ,  0 , None , !�F Index , Arial ,  10 ,  180 ,  250 ,  20�    60 ,  0 ,  0 ,  0 , None , !�I Glossary , Arial ,  10 ,  1�    , None , !�I Glossary , Arial ,  10 ,  180 ,  250 ,  20 , �   abel , Arial ,  12 ,  180 ,  250 ,  20 ,  60 ,  0 , -1 ,  0�   0 ,  20 ,  60 ,  0 , -1 ,  0 , None , !�V Glossary Letter L�   None , !�V Glossary Letter Label , Arial ,  12 ,  180 ,  25�   l , Arial ,  12 ,  180 ,  250 ,  20 ,  60 ,  0 , -1 ,  0 , �     20 ,  60 ,  0 , -1 ,  0 , None , !�V Glossary Letter Labe�   e , !�V Glossary Letter Label , Arial ,  12 ,  180 ,  250 ,�    Arial ,  12 ,  180 ,  250 ,  20 ,  60 ,  0 , -1 ,  0 , Non�   0 ,  60 ,  0 ,  0 ,  0 , None , !�V Glossary Letter Label ,�    0 ,  0 , None , !�F Index , Arial ,  10 ,  180 ,  250 ,  2�   , !�F Index , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 , �   rial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None �   80 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�F Index , A�    ,  60 ,  0 ,  0 ,  0 , None , !�F Index , Arial ,  10 ,  1�   80 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�I Glossary �   ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�D Bar ,�    ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�D Bar , Arial ,  10 �   ,  0 ,  0 ,  0 , None , !�D Bar , Arial ,  10 ,  180 ,  250�   0 , None , !�D Bar , Arial ,  10 ,  180 ,  250 ,  20 ,  60 �   D Bar , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  �    ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !��     250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�F Image , Arial�   60 ,  0 ,  0 ,  0 , None , !�F Image , Arial ,  10 ,  180 ,�    0 , None , !�F Image , Arial ,  10 ,  180 ,  250 ,  20 ,  �    Image , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 , �   ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�F�    250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�F Image , Arial �     0 ,  0 ,  0 , None , !�I Glossary , Arial ,  10 ,  180 , �   ne , !�I Glossary , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,�   , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , Noj�    Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , Non�   ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,�   1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  �   e , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !��   !�;  , Arial ,  10 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 , Non�    ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , �   0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0�    0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  �   ,  0 ,  0 ,  0 , None , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 , �    ,  0 ,  0 , None , !�;  , Arial ,  10 ,  0 ,  0 ,  0 ,  0 �   ne , !�F Table , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0�   , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , No�     180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�F Table �    20 ,  60 ,  0 ,  0 ,  0 , None , !�F Table , Arial ,  10 ,�   ,  0 ,  0 , None , !�F Table , Arial ,  10 ,  180 ,  250 , �   e , !�F Table , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 "�     0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�;  , Arial ,  10 ,�    0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 , None , !�1  ,  ,  0 ,  0�    0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�;  , Arial ,  10 , �     0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 , �     ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,�    , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1�   �;  , Arial ,  10 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 , None�   ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�    ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 �   0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0�     0 ,  0 ,  0 , None , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  �     0 ,  0 ,  0 ,  , !�;  , Arial ,  10 ,  0 ,  0 ,  0 ,  0 ,�   ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,�    ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 �   0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0�     0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 , None , !�1  ,  ,  0 ,  ��    ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 �    oder weniger vollst�ndige Aufzeichnungen gibt, die aber, d�   spekt war, da� es an verschiedenen Stellen im Internet mehr�   ationen vielleicht f�r immer verloren gehen. Ein weiterer A�   eitung und �berblick!�
 /N /Just L!�/P /Just L /Text Ursp�   r�nglich war dieses Programm nur dazu gedacht, die INVISICL�   UES(TM) zu den alten INFOCOM-Adventures in elektronischer F�   orm wiederaufzubereiten, um zu verhindern, da� diese Informm  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�   st neu in Version 1.1 ?!�F /L /Jump Referenzen /Link /Macro�   as ist neu... /Link /Macro /Play /popup /Just L /Text Was i�   192,192), 0!�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  9   �% /H /Just L /Text The Hint Library 1.1!�$ /T /Just L /Tex     0 ,  0 ,  0 ,  , !�                                       �     0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 , �   ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,   a normalerweise nur als Textdatei verf�gbar, der eigentlich  e zur Verf�gung zu stellen (und nicht nur unbedingt f�r Com�    aufgefordert, anderen Leuten seine besten Tips und Hinweis�   , eine Hinweis-Bibliothek aufzubauen und jeder wird hiermit�   ssammlungen anzulegen. Das nunmehr verfolgte Ziel soll sein�   ignet ist, sondern auch die M�glichkeit bietet, neue Hinwei�   ger�ckt, das nicht nur zum Lesen solcher Hinweisdateien gee�   nn immer mehr der Gedanke an ein System in den Vordergrund �   nehmen will.����Bei der Entwicklung dieses Programms ist da�   nd man selber dosieren kann, wieviel Hilfe man in Anspruch �   ich raubt, indem man in einer Komplettl�sung zuviel sieht u�   sammlungen ist, da� man sich den Spielspa� nicht versehentl�   de) Hinweise zu geben. Der gro�e Vorteil an solchen Hinweis�   blemstellen in den Textadventures (in der Pr�zision steigen�   Idee hinter den InvisiClues(tm) war es zu verschiedenen Pro�   en Idee dieser Hinweissammlungen nicht gerecht werden. Die �  puterspiele !). Um f�r m�glichst viele Menschen dieses Prog  t ausw�hlen. Das versehentliche Lesen von Hinweisen soll ni  en Sie Informationen nur lesen k�nnen, wenn Sie sie explizi  e zur Verf�gung stehenden Hinweise zum Lesen an. Dabei werd  eser bietet Ihnen, normalerweise nach Themen gegliedert, di  Teilen.  Da ist zum einen der Reader, der "Lese"-Teil. Di  zum Programm selber:��Es besteht im  wesentlichen aus zwei   inen Umst�nden kommerziell genutzt werden darf.����Und nun   lich dem Sammeln von Informationen dienen soll und unter ke	   soll hier nochmal betont werden, da� das System ausschlie�
  te, damit wir das weitere Vorgehen besprechen k�nnen.����Es  usammenzustellen. In diesem Falle kontaktieren Sie mich bit  erkl�ren w�rde, ein weiteres Sprachpaket f�r das Programm z  n. Ich w�rde mich also sehr freuen, wenn sich jemand bereit  n von der Oberfl�che und der Online-Hilfe unterst�tzt werde  ramm nutzbar zu machen, sollen auch m�glichst viele Sprache   cht m�glich sein. Zur Zeit begegnen Ihnen im Reader folgend!    PCX-,TGA- und JPEG-Dateien verwendet. Zu erreichen unter:  eile seines MPICVIEW-Projekt werden von mir zur Anzeige von  Personen gilt mein besonderer Dank:����Detlef Meister. T  '  G��� 
� - 4 M     � Topic@Einleitung  �      �  	  � 2000   �  ��;�   =  �8 Sprachdateien;Sprachen;  Hinweisdateien;Infocom;�berblick;�� F�     �
 Einleitung�   �� U�     �  �� 	�  U-�   !�) /T /Just L /Text Einl  �    �    �  ��;�   1  �, Autor;Borland Delphi;Inform  ation;Danksagung;�� B�     �
 Referenzen�� Q�     �    �� 	��  �-�   !� /T /Just L /Text Referenzen!�
 /N /Ju  st L!��/P /Just L /Text Autor: Stefan Meier����Folgenden �  rtrag /Link /Macro /Play /popup /Just L /Text Lizenzbedingu   /Play /popup /Just L /Text Referenzen!�P /L /Jump Lizenzvew  MIDI, AVI,...)��Weiteres finden Sie unter Hinweis-Dateien-l  e��Hinweistypen: Texte, Bilder und Multimediadateien( z.B. j0  ��Meister@rz.fhtw-berlin.de����Allen Ex-Infocomlern, die mi#  migung entbindet den H�ndler nicht von den anderen Pflichte$  n, die sich aus diesem Vertrag ergeben.����Mein besonderer %  Dank gilt Detlef Meister f�r sein Freeware-Projekt MPICVIEW&  .��Dieses Programm nutzt Teile dieses Projektes zum Anzeige'  n von JPEG, TARGA und PCX-Dateien.��Sie erreichen Detlef Me(  ister unter;��Meister@rz.fhtw-berlin.de�� ��Kontaktadresse)  :��Stefan Meier, Erfstr. 65, D-52249 Eschweiler, Germany��*  AOL:��SMeier7777��E-Mail:��SMeier7777@aol.com��Stefan.M    eier@post.rwth-aachen.de  
� �                               �                                                          �  	  � 1000   �  ��7i     � �berblick;Inhalt;�� B�     �  �n�� 
� - 4 I     � Topic@Referenzen  �        twickelt.��  
� �                                        .  .������The Hint Library 1.1 wurde mit Borland Delphi 2.0 en/  t Ihren Textadventures Computergeschichte geschrieben haben""   des Programms aufh�ren.��Das Widerrufen der Vertriebsgeneh3   einer besonderen schriftlichen Genehmigung.��Kein H�ndler 4  darf mehr als 12 DM (oder den entsprechenden Betrag in ande5  ren W�hrungen, z.B. $8 US) f�r die Verbreitung dieses Progr6  amms verlangen.����Alle THL-Dateien eines H�ndlers m�ssen a7  uf eine m�glichst kleine Menge Disketten verteilt werden. D8  ie Verteilung mittels einer unnat�rlich gro�en Menge Disket9  ten ist VERBOTEN.��F�r solche Disketten, auf denen THL-Date:  ien vertrieben werden, d�rfen unter keinen Umst�nden mehr a;  ls 12 DM (oder der entsprechende Betrag in anderen W�hrunge<  n, z.B. $8 US) verlangt werden.��Diese Bedingungen gelten s=  owohl f�r die Verbreitung dieses Programms, als auch f�r al>  le THL-Dateien, die von anderen Autoren erstellt werden.���?  �Die Genehmigung zur Verteilung des Programms kann schriftl@  ich widerrufen werden. Sp�testens 30 tage nach dem Ausstell1  ungsdatum des Widerrufs, mu� der H�ndler mit der Verteilung�2  der Verbreitung �ber "Magazin-CDs" oder "Magazin-Disketten"C  , die aus der direkten oder indirekten Nutzung des ProgrammD  s entstehen, auch dann nicht, wenn der Autor auf m�gliche SE  ch�den durch die Nutzung des Programmes hingewiesen worden F  ist. ����Wenn Sie beabsichtigen, mit dem Programm THL-DateiG  en zu erstellen und zu verbreiten. sollten Sie mir mitteileH  n, welches Projekt sie vorhaben und zuerst bei mir anfragenI  , ob jemand anders gerade an einem THL-File zu dem jeweiligJ  en Thema schreibt. Obwohl das Programm unentgeldlich benutzK  t werden darf, ist es unter KEINEN UMST�NDEN ERLAUBT, f�r "L  eigene" THL-Files in irgendeiner Form Geb�hren zu verlangenM  . Wenn Sie Ihre THL-Dateien zur Verf�gung stellen wollen, sN  ollten Sie mir eine Kopie zukommen lassen. Der einfachste WO  eg ist, die Datei an der unten angegebenen FTP-Adresse abzuP  legen. �� ��Die Verbreitung �ber Warenh�user bedarf einer bA  esonderen schriftlichen Genehmigung.��Ebenso bedarf es bei �B  Stefan Meier, tr�gt in keinem Falle die Haftung f�r Sch�denS  n und m�ssen alle Kopien davon l�schen.��Dieses urheberrechT  tllich gesch�tzte Programm wird als "Freeware" vertrieben. U  Sie d�rfen das Programm unentgeldlich benutzen und an anderV  e weitergeben.��Alle Rechte an diesem Programm geh�ren StefW  an Meier und werden durch das Urheberechtsgesetz der BundesX  republik Deutschland und internationale��Abkommen gesch�tztY  . Daher mu� das Programm wie anderes gesch�tztes Material bZ  ehandelt werden (z.B. B�cher und Tontr�ger).����Dieses Prog[  ramm darf nicht vermietet werden. Au�erdem ist es nicht erl\  aubt, das Programmpaket zu ver�ndern, zu �bersetzen, zu dis]  sassemblieren oder zu decompilieren.��Wenn Sie eine der Bed^  ingungen dieses Vertrages verletzen, erlischt automatisch I_  hr Nutzungsrecht f�r dieses Programm und Sie m�ssen alle Ko`  pien l�schen.����Das Programm und die Dokumentation werden Q  so zur Verf�gung gestellt, "wie sie sind", d.h. der Autor, R  t einverstanden sind, d�rfen Sie das Programm nicht benutzeq  11\HELPFILE\DATEIM~1.BMP /Just L /Text Mit Datei �ffnen wb  t L /Text Die Programm-Men�s:!�8/R /Link E:\WORK\HINT_R~1.c  t L /Text Hiermit beenden Sie The Hint Library!�& /H 2 /Jusd  nden!�a /R /Link E:\WORK\HINT_R~1.11\HELPFILE\EXIT.BMP /Juse  ie unter anderem die Programmversion und Kontaktadressen fif   /Just L /Text Hiermit �ffnen Sie ein Infofenster, in dem Sg  atei auf.!�� /R /Link E:\WORK\HINT_R~1.11\HELPFILE\INFO.BMPh  P.BMP /Just L /Text Mit diesem Knopf rufen Sie diese Hilfedi  ie den Editor.!�m /R /Link E:\WORK\HINT_R~1.11\HELPFILE\HELj  R~1.11\HELPFILE\EXISTF~1.BMP /Just L /Text Hiermit �ffnen S�   Editor-Eintr�gen via Drag & Drop��Erweitertes Save/Compile�   !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�o  enzvertrag!�
 /N /Just L!��/P /Just L /Text Bitte lesen Sip  e diesen Lizenzvertrag komplett bevor Sie dieses Programm ba  enutzen. Wenn Sie mit den Bedingungen dieses Vertrages nich��  �hlen Sie eine Hinweissammlung aus und �ffnen den "Reader"��  ich bitte, um das weitere Vorgehen abzusprechen. ��Mit Sprr  rf�gung stellen k�nnten. In diesem Falle kontaktieren Sie ms  r dar�ber freuen, wenn Sie mir ein neues Sprachpaket zur Vet  uen Sie bitte auf der THL-Homepage nach. Ich w�rde mich sehu  diesem Programm hinzugef�gt werden.F�r andere Sprachen schav  chpaket mitgeliefert. Zus�tzliche Pakete k�nnen einfach zu w  n. Standardm��ig wird mit diesem Programm das deutsche Sprax  ie einen Dialog, in dem Sie ein Sprachpaket ausw�hlen k�nney  1.BMP /Just L /Text Mit Sprache - Sprache w�hlen �ffnen Sz   Formular.!��/R /Link E:\WORK\HINT_R~1.11\HELPFILE\SPRACH~{   Mit Editor �ffnen Sie das Editorfenster mit einem leeren|  ink E:\WORK\HINT_R~1.11\HELPFILE\EDITOR~1.BMP /Just L /Text}  der.��Mit Beenden verlassen Sie The Hint Library!�� /R /L~  ammlung nach ihrem behandelten Titel aus und �ffnen den Rea  �Mit Datei �ffnen (�ber Titel)... w�hlen Sie ein Hinweiss"�  acheinstellung speichern k�nnen Sie bestimmen, ob die eing�  um Umgang mit dem Windows Hilfesystem��Info zeigt Ihnen e�  T_R~1.11\HELPFILE\OPENBTN.BMP /Just L /Text Hiermit �ffnen �  Sie eine THL-Datei zum "Hinweis-Lesen". Hinweise zum Umgang�   mit dem Reader finden Sie unter THL-Hinweis-Dateien lesen!�  �� /R /Link E:\WORK\HINT_R~1.11\HELPFILE\VOPEN.BMP /Just L �  /Text Auch hiermit k�nnen Sie eine THL-Datei zum Lesen �ffn�  en, allerdings sehen Sie hier nicht die Dateinamen, sondernk   die Titel der Hinweissammlungen.!�_ /R /Link E:\WORK\HINT_�  lw�rtern suchen��Hilfe-benutzen zeigt Ihnen Erkl�rungen z�  - Suchen k�nnen Sie in der ganzen Hilfedatei nach Schl�sse�  lfedatei auf und starten im Inhaltsverzeichnis��Mit Hilfe �  1.BMP /Just L /Text Mit Hilfe - Inhalt rufen Sie diese Hi�  aden wird.!��/R /Link E:\WORK\HINT_R~1.11\HELPFILE\HILFEM~�     � Inhaltsverzeichnis�� Q�     �  �� 	rh  �-�   !�  estellte Sprache beim n�chsten Start automatisch wieder gel"�  in Fenster, dem Sie die aktuelle Programmversion, Kontaktad�    �  �� 	�h  �-�   !�  /T /Just L /Text Wo gibt es... �  teien;Neue Versionen;�� I�     � Wo gibt es ?�� X�   �    �  	  � 8000   �  ��>�   .  �) Sprachdateien;THL-Da�  q  /[�� 
� 0 7 P     � Topic@Wo gibt es...  �  �   /Just L!�t /L /Jump Was sind THL Dateien... /Link /Macro /�  �� 	�P  �-�   !� /T /Just L /Text Der THL-Editor!�
 /N�  ateien,editieren;�� F�     �
 Der Editor�� U�     �  �  �  	  � 5000   �  ��;�   -  �( THL-Editor;Editor;THL-D�  wahlliste unten k�nnen Sie direkt zu verwandten Themen spri  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !� �  �   a�� 
� 6 = V     � Topic@Das Hinweis FensterI    �=�� 
 = D ]   %  �  Topic@Das Hinweis Editierfe�  >  ֮�� 
{ : A Z   "  � Topic@Das Bildanzeige Fenst�  , Bedienung;Editor;�� U%    � Die Bedienung des Editor    ressen und weitere Informationen entnehmen k�nnen  
� �  �  %  �Z�� 
� : A V   "  � Topic@Was sind THL Dateien.�  en.��Wenn Sie eigene Dateien entwerfen, verwahren Sie immer�  G: THL-Dateien k�nnen nicht mehr im Editor bearbeitet werd�  en gespeichert, allerdings ohne sie zu �bersetzen.��ACHTUN�   SEHR EMPFOHLEN !). In einer THR-Datei werden die Editordat�  /B /Just L /Text Ggf. Abspeichern der Daten als THR-Datei (�  r Hinweise und Benennen von Bildern u.�. mit dem Editor!�D�  teien verl�uft wie folgt:!�U /B /Just L /Text Eingeben alle�   dieses Programms.��Die prinzipielle Entstehung von THL-Da�  ht mit einem Texteditor lesbar, sondern nur mit dem Reader�  der und Multimediadateien enthalten. Diese Dateien sind nic�  P /Just L /Text THL-Dateien sind Bin�rfiles, die Texte, Bil�  2-�   !� /T /Just L /Text THL-Dateien!�
 /N /Just L!�/�  �     � Was sind THL Dateien...�� ^�     �  �� 	�  �  eien;Hinweise;Bilder;Formate;THL-Dateien;THR-Dateien;�� O�  ..  �    �    �    �  ��H�   H  �C Multimedia-Dat��   eine Kopie der THR-Datei !!!!�= /B /Just L /Text �bersetze�  Play /popup /Just L /Text Was sind THL-Dateien und wie ents�  er, da� jeder diese Hinweise lesen/ansehen/h�ren kann.  
��  re Formate unterst�tzt, allerdings ist dann nicht mehr sich�  t werden WAV, AVI, MIDI, MOV. Prinzipiell werden auch weite�  ersehen.!�� /B /Just L /Text Multimedia-Dateien, unterst�tz�  s Bildern definieren und diese mit eigenen Beschreibungen v�  ga��Besonderheiten: Sie k�nnen mit dem Editor Auschnitte au�   /Text Bilder, unterst�tzte Formate: Bitmap, JPeg, PCX, Tar�   /Just L /Text Texte ( ein- oder mehrzeilig )!�� /B /Just L�  mehr enthalten. Folgende Typen von Hinweisen gibt es:!�/ /B�  se enthalten, allerdings k�nnen Hinweise keine Unterthemen �  erschiedene Themen. Ein Thema kannn Unterthemen oder Hinwei�   /Just L /Text Normalerweise enth�lt eine Hinweissammlung v�  �2 /H 1 /Just L /Text Der Aufbau von THR/THL-Dateien:!�� /P�  n der Editordaten in eine THL-Datei!� /H 1 /Just L /Text !�  tehen sie?!�| /L /Jump Eigenentwicklung von Hinweissammlung�  klaren, fragen Sie beim Inhaber der Urheberrechte um Erlaub�  nis.!�1/B /Just L /Text Verbreiten sollten Sie normalerwei�  se nur die THL-Datei, damit au�er Ihnen keine die Daten ver�  �ndern kann. WICHTIG: Behalten Sie aber immer eine Kopie �  der THR-Datei, da sie sonst auch selber Ihre Daten nicht me�  hr �ndern k�nnen. EINE THL-DATEI KANN NICHT MEHR IM EDITOR �  VER�NDERT WERDEN !!�E/B /Just L /Text Lassen Sie mir eine �  Kopie Ihrer THL-Datei zukommen. Am einfachsten geht dies, i�  p://members.aol.com/thlhome/incoming��Sie k�nnen mir auch �  eine Diskette per Post schicken, oder mir eine Adresse im I+  nternet benennen, unter der die Datei erh�ltlich ist  
� �  ndem Sie die Datei an die folgende ftp-Adresse senden:��ft�  Y  ��� 
� - 4 M     � Topic@Der Editor  �    4  eigener THL-Dateien.!�d /L /Jump Die Bedienung des Editors �  en /Link /Macro /Play /popup /Just L /Text Die Entwicklung j�  Form zu �bertragen. Sind Sie sich �ber die Rechtslage im un�   sollten Sie folgende Hinweise beherzigen:!�d/B /Just L /T�  ext Bevor Sie mit Ihrer Arbeit beginnen, kontaktieren Sie m�  ich, um zu erfragen, ob schon jemand anderes an einer Datei�   zu Ihrem Spiel / Thema arbeitet. Dies soll einerseits verh�  indern, da� Arbeit unn�tigerweise doppelt gemacht wird und �  andererseits gibt es mir die M�glichkeit, einen �berblick ��  ber die Entwicklung des THL-Projekts zu bewahren!�� /B /Jus�  t L /Text �berlegen Sie sich eine Gliederung f�r Ihre Hinwe�  issammlung. Wo treten Fragen auf ? Wo kann man Sinnabschnit�  te abgrenzen? Wo ist Bildmaterial hilfreich ?!�� /B /Just L�   /Text Vergleichen Sie Ihre L�sungswege, wenn m�glich, mit �  anderen L�sungen, um Fehler oder Auslassungen zu vermeiden.�  !�'/B /Just L /Text Bitte achten Sie darauf, da� Sie keine�   Urheberrechte verletzen. So ist es normalerweise nicht erl�  aubt, kommerziell vertriebene "Hintbooks" in elektronische ��  n, eigene Hinweissammlungen zu entwerfen und zu verbreiten,    s.aol.com/smeier7777/thlfiles  
� �                     �  aol.com/smeier7777/thl_lang����THL Dateien:��ftp://member�  .aol.com/tinyyeti/thl1.d����Sprachpakete:��ftp://members.�  ie FTP Zugriff bevorzugen:����THL Software:��ftp://members�  mbers.aol.com/thlhome/index.htm!�� /B /Just L /Text Wenn S�   Sprachpakete und THL-Dateien findet man unter:��http://me`    !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  ngen!�> /P /Just L /Text ������The Hint Library � 1996-97 S�    �  	  � 7000   �  ��>�   8  �3 Benutzung, Bedingung�  en;Vertriebsbedingungen;Lizenz;�� I�     � Lizenzvertran  g�� X�     �  �� 	��  
-�   !� /T /Just L /Text Liz�   Entwicklung;Eigene Dateien;THL-Dateien;�� ^�   +  �& Eig�  enentwicklung von Hinweissammlungen�� m�     �  �� 	��    -�  	 !�0 /T /Just L /Text Entwicklung eigener THL-Date�  ien!�
 /N /Just L!�� /P /Just L /Text Wenn Sie beabsichtige"�  *  �2�� 
� 1 8 Q     � Topic@Der THL Reader  �    elwort PIC und Multimediadateien MM. Bei Themen sehen Sie s�  or ihrem Eintrag das Schl�sselwort HINT, Bilder das Schl�ss�  sehen Sie Ihr Projekt als Baumansicht, Hinweise enthalten v�  E ZUM ERSTELLEN VON THL-DATEIEN !!��/E /Just L /Text Hier �   /Just L!�P /P /Just L /Text BITTE BEACHTEN SIE DIE HINWEIS�  -Men���Sicherheitsabfrage beim Schlie�en des Editors  
� �  Hinweissammlungen  �    �    �    �  ��W�   ,  �'�  E:\WORK\HINT_R~1.11\HELPFILE\EDITOR.BMP /Macro /Play /Popup�   Bedienung des THL-Editors!�
 /N /Just L!�R /I /Jump /Link �  s�� d5    �  �� 	�  t-�   !�. /T /Just L /Text Die�  /Just L /Text Bedeutung der Kn�pfe:!�� /R /Link E:\WORK\HIN�    �  	  � 4000   �  ��?�   &  �! Hinweise lesen;THL-    ngen.  
� �                                                  tefan Meier  
� �                                            �  !�  !�                                                  "  ie ersten Buchstaben des Titels. Wenn Sie neue Eintr�ge hin  a� z.B. Video-Dateien in der Regel relativ gro� sind und de  edia-Editierfenster ge�ffnet. Bitte beachten sie hierbei, d  Dateien zu Ihrem Projekt hinzuzuf�gen. Dazu wird das Multim   /Just L /Text Knopf Nummer 5 erlaubt es Ihnen, Multimedia-  f�gen. Dazu wird das Hinweis-Editierfenster ge�ffnet.!��/E  sem Knopf k�nnen Sie einen neuen Hinweis in Ihr Projekt ein  Bildbereiche definieren k�nnen.!�� /E /Just L /Text Mit die  n neuen Bildeintrag zu Ihrem Projekt hinzuf�gen k�nnen und 	  t Hier �ffnen Sie das Bild-Editierfenster, mit dem Sie eine
  wird das Themen-Editierfenster ge�ffnet.!�� /E /Just L /Tex  k�nnen Sie Ihrem Projekt ein neues Thema hinzuf�gen. Dabei   gen k�nnen.!�� /E /Just L /Text Bei Dr�cken dieses Knopfes   n�pfe 2-5 je nachdem, was Sie f�r diesen Eintrag noch einf�  zer". Wenn Sie ein Element selektieren ver�ndern sich die K  zuf�gen, fungiert der jeweis selektierte Eintrag als "Besit   mentsprechend Ihre THL-Datei anw�chst. Obwohl die Multimedi!   M�glichkeit einen Eintrag innerhalb seiner Ebene nach oben  machen usw.!�� /E /Just L /Text Dieser Knopf gibt Ihnen die  ndern, d.h. Sie k�nnen nicht aus einem Thema einen Hinweis   �ffnet. Es ist nicht m�glich den Typ eines Eintrags zu ver�  ndern. Je nach Typ wird das entsprechende Editierfenster ge  t Mit diesem Knopf k�nnen Sie den selektierten Eintrag ver�  r Beschreibung des Verkn�pfungsfensters.!�/E /Just L /Tex  zu anderen Eintr�gen definieren. Weiteres finden Sie bei de   k�nnen Sie zum aktuell selektierten Eintrag Verkn�pfungen   eader nicht versteckt dargestellt.!�� /E /Just L /Text Hier  Information in Ihr Projekt einf�gen. Diese wird sp�ter im R  !�� /E /Just L /Text Mit diesem Knopf k�nnen Sie eine neue   dia-Formate u.U. f�r manche Benutzer nicht mehr lesbar sind  bh�ngen, sollten Sie daran denken, da� ausgefallene Multime  a-Unterst�tzung alleine von den F�higkeiten Ihres Systems a�0   zu verschieben. Auch wird werden evt. vorhandene Untereint1  r Schriftarten verwenden, die beim System mitgeliefert werd"   sind. Um unerw�nschte Effekte zu vermeiden, sollten Sie nu#  arten zur Verf�gung haben, die auf Ihrem System installiert$  te beachten Sie, da� andere Benutzer evt.nicht alle Schrift%  ie im Reader benutzt wird, um Ihren Titel darzustellen. Bit&   Mit dem Schrift-Knopf k�nnen Sie eine Schriftart w�hlen, d'  amit Ihr Projekt �bersetzt werden kann.!�u/E /Just L /Text(  ter im Reader erscheint. Dieses Feld mu� ausgef�llt sein, d)  ekt an. Dies ist kein Dateiname, sondern der Titel, der sp�*  ust L /Text In diesem Feld geben Sie den Titel f�r Ihr Proj+   Sie vorsichtig bei der Benutzung dieser Funktion.!�� /E /J,  ventuell vorhandene Untereintr�ge werden mitgel�scht. Seien-  f l�schen Sie den momentan selektierten Eintrag. Achtung: E.  Verschieben nach unten"!�� /E /Just L /Text Mit diesem Knop/  r�ge mit verschoben!�; /E /Just L /Text Analog zu Knopf 9 "�@  en.!�� /E /Just L /Text In diesem Feld geben Sie Informatio3  mas ein. Schlie�en Sie das Fenster mit OK, wird das Thema z    u Ihrem Projekt hinzugef�gt.  
� �                       �  /Link /Macro /Play /popup /Just L /Text Die Bedienung des Ez  et sich ein Popup-Men�, mit dem Sie direkt neue Eintr�ge er5  n Sie in der Baumansicht die rechte Maustaste dr�cken, �ffn6   /Just L /Text Sonstige Funktionen:!�4/P /Just L /Text Wen7  �nnen Sie Ihr Projekt in eine THL-Datei �bersetzen.!�' /H 18  ichern und den Editor verlassen.��Mit dem Compiler-Men� k9  it dem Datei-Men� k�nnen Sie Ihre Datei im THR-Format spe:  eben!� /H 1 /Just L /Text Die Men�s:!�� /P /Just L /Text M;  lichkeit, zus�tzliche Informationen zu Ihrem Projekt einzug<  Hummel.!�n /E /Just L /Text Dieses Feld gibt Ihnen die M�g=  Written 1997 by Harry Hummel oder Copyright � 1997 Harry >   sein, damit das Projekt �bersetzt werden kann. Beispiel: ?  nen �ber sich als Autor an. Auch dieses Feld mu� ausgef�llt2   /P /Just L /Text Unter Text tragen Sie den Titel Ihres The�  r Hinweis zum aktuell selektierten Thema hinzugef�gt.  
� B  Hinweis ein. Wenn Sie das Fenster mit OK schlie�en, wird deC  up /Just L!�� /P /Just L /Text Unter Text tragen Sie Ihren D  E:\WORK\HINT_R~1.11\HELPFILE\HINTEDIT.BMP /Macro /Play /PopE  Das Hinweis-Editierfenster!�
 /N /Just L!�T /I /Jump /Link F  ster�� e�     �  �� 	�	  <-�   !�+ /T /Just L /Text G  eingabe;Text;Hinweis;�� V�     � Das Hinweis EditierfenH  nster  �    �  	  � 5020   �  ��K�   !  � HinweisK  �  R��� 
� < C \   $  � Topic@Das Themen EditierfenL  ster  �    �  	  � 5030   �  ��J~     � ThemeneiM  ngabe;Text;�� U�     � Das Themen Editierfenster�� d�N       �  �� 	��  .-�   !�* /T /Just L /Text Das Themen-P  Editierfenster!�
 /N /Just L!�S /I /Jump /Link E:\WORK\HINT_  r>!�1 Bild-Editierfenster,Das Bilder Editierfenster, 0,!�' A  _R~1.11\HELPFILE\TOPEDIT.BMP /Macro /Play /Popup /Just L!���  .11\HELPFILE\MAIN.BMP /Just L!� /H /Just L /Text !�( /H 2 a  eschreibung hinzuf�gen. Wenn Sie eine neue Datei ausw�hlen,R  hrer Bereichsliste hinzugef�gt. Sie m�ssen dann noch eine BS  ald Sie die linke Maustaste loslassen, wird der Auschnitt IT  d markieren den Bildauschnitt, den Sie benennen wollen. SobU  ustaste in das Bild, halten die linke Maustaste gedr�ckt unV   Bildhinweise eintragen. Dazu klicken Sie mit der linken MaW  ichseditor k�nnen Sie separate Bildausschnitte als einzelneX  wird die jeweils behandelte Bilddatei eingetragen.  Im BereY  Macro /Play /Popup /Just L!�:/P /Just L /Text Unter Datei Z  S /I /Jump /Link E:\WORK\HINT_R~1.11\HELPFILE\PICEDIT.BMP /[   /T /Just L /Text Das Bilder-Editierfenster!�
 /N /Just L!�\   Bilder Editierfenster�� d�     �  �� 	��  �-�   !�*]  ten;Bilder;Fortschrittsanzeige;Bereiche;�� U�     � Dash  Der THL-Editor,(Global), 0,<Der Editor>!�' Der-THL-Editor,(�  �  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  p   wird automatisch das komplette Bild als Bereich eingetragec   /Just L /Text Das Multimedia-Editierfenster!�
 /N /Just L!d  �R /I /Jump /Link E:\WORK\HINT_R~1.11\HELPFILE\MMEDIT.BMP /e  Macro /Play /Popup /Just L!�� /P /Just L /Text Unter Datei f  tragen Sie die behandelte Multimedia-Datei ein. Unter Beschg  reibung geben Sie der Datei einen Titel. Wenn Sie das Fenst�  er mit OK schlie�en, wird dieser Multimedia-Eintrag zum akt}  Global), 0,<Der Editor>!�Q Eigene THL-Dateien erstellen,(Gl�   zu diesem Bild definieren, wird immer der erste Bereich (ni  nzelner Hinweis behandelt.��WICHTIG: Wenn Sie Verkn�pfungenj  wird sp�ter im Reader jeder eingetragene Bereich als ein eik  Obwohl Sie im Editor nur einen Eintrag f�r ein Bild sehen, l  ag zu dem aktuell selektierten Thema hinzugef�gt. Beachte: m  . Wenn Sie das Fenster mit OK schlie�en, wird der Bildeintrn  ie diesen eintrag nicht w�nschen, ihn aus der Liste l�scheno  n. Sie sollten die Beschreibung hierzu �ndern, oder falls S"b  edia Editierfenster�� h�     �  �� 	�c  �-�   !�. /T�  itor und zum Erstellen von THL-Dateien finden Sie unter Derr  PEG, TARGA, PCX) in Ihre Dateien aufnehmen.��N�heres zum Eds  Sie Multimediadateien ( Sound, Videos ) und Bilder ( BMP, Jt  komfortabel in einem Fenster erledigt. Neben Texten k�nnen u  ichkeit gibt, neue Hinweis- Dateien anzulegen. Dieses wird v  esen.��Der andere Teil ist der Editor, der Ihnen die M�gl�  >!�5 Hinweis-Editierfenster,Das Hinweis Editierfenster, 0,!x  nweis Fenster>!�* Hinweis-Dateien-lesen,(Global), 0,<(None)�  zeugen k�nnen.��Zus�tzlich k�nnen Sie Eintr�ge innerhalb dey  issammlungen>!�8 Hinweis-Anzeigefenster,(Global), 0,<Das Hi{  LEN VON THL-DATEIEN,(Global), 0,<Eigenentwicklung von Hinwe|  obal), 0,<Eigenentwicklung von Hinweissammlungen>!�N ERSTEL  l  R��� 
� @ G `   (  �# Topic@Das Multimedia Editie�  rfenster  �    �  	  � 5040   �  ��N�   *  �% Multq  imedia-Dateien;Dateibeschreibung;�� Y�   "  � Das Multim��  -THL-Editor. ( Bitte unbedingt lesen ! )��Nicht zu sehen is�   wird eine Warnung erscheinen, wenn Sie beispielsweise Hinw�  ��Da die Hinweise einer Auswahl in der Pr�zision ansteigen,�  nw�hlen, �ffnet sich das Hinweis-Anzeigefenster. Anmerkung:�   F�r Hinweise. Wenn Sie durch Doppelklicken einen Hinweis a�  Link E:\WORK\HINT_R~1.11\HELPFILE\HINTPIC.BMP /Just L /Text�  n oder Hinweise. Diese sehen in etwa wie folgt aus:!�l/R /�  e eine Ebene tiefer. Dort finden Sie entweder weitere Theme�  enth�lt. Durch doppeltes Anklicken eines Themas gelangen Si�  r in der mitte sehen Sie die Hauptthemen, welche die datei �  /Popup /Just L!�/P /Just L /Text In dem Aufz�hlungsfenste�  /Link E:\WORK\HINT_R~1.11\HELPFILE\READER.BMP /Macro /Play �  n einer THL-Datei sehen Sie folgendes Fenster:!�R /I /Jump �  N /Just L!�\ /P /Just L /Text Nach der �ffnen und �bersetze�   �� 	�!  g-�  	 !� /T /Just L /Text Der THL-Reader!�
 /�  Reader;Reader;�� J�     � Der THL Reader�� Y�     � ��  eis 3 lesen wollen, bevor Sie die Hinweise 1 und 2 gelesen �  Kontrolle;Multimediadateien abspielen;Multimediaplayer;�� �  r  �    �  	  � 4030   �  ��G�   G  �B Multimedia-�  �5 Informationsfenster,(Global), 0,<Informationsfenster>!�Z�  eis-Fenster!�
 /N /Just L!�T /I /Jump /Link E:\WORK\HINT_R~�  ^�     �  �� 	��  �-�   !�$ /T /Just L /Text Das Hinw�  weis;Hinweis zeigen;�� O�     � Das Hinweis Fenster�� �    �    �  	  � 4020   �  ��D�   '  �" Verdeckter Hin�  C.BMP /Just L /Text F�r Informationen. Durch einen Doppelcl�  igefenster.!�� /R /Link E:\WORK\HINT_R~1.11\HELPFILE\INFOPI�   Doppelklicken ein Bild anw�hlen, �ffnet sich das Bild-Anze�  ELPFILE\PICPIC.BMP /Just L /Text F�r Bilder. Wenn Sie durch�  ltimedia-Kontrollfenster.!�� /R /Link E:\WORK\HINT_R~1.11\H�  klicken eine Multimedia-Datei ausw�hlen, �ffnet sich das Mu�  Just L /Text F�r Multimedia-Hinweise. Wenn Sie durch Doppel�  haben.!�� /R /Link E:\WORK\HINT_R~1.11\HELPFILE\MMPIC.BMP /��  R�     � Das Multimedia Fenster�� a�     �  �� 	�� �  eis innerhalb der momentan g�ltigen Auswahlliste als Gelese�  t  "Schlie�en" das Fenster zumachen. Dabei wird dieser Hinw�  ie den Knopf "Hinweis zeigen" dr�cken. Danach k�nnen Sie mi�  hen Sie das folgende Fenster. Um den Text zu lesen, m��en S�  P /Just L /Text Wenn Sie einen Hinweis ausgew�hlt haben, se�  1.11\HELPFILE\HINTVIEW.BMP /Macro /Play /Popup /Just L!�,/�  ,<Das Multimedia Editierfenster>!�? Multimedia-Kontrollfens�   Multimedia-Editierfenster,Das Multimedia Editierfenster, 0�  e Abspielvorg�nge werden automatisch gestoppt. �ber die Aus�  �nnen. Mit OK schlie�en Sie das Fenster. Dabei noch laufend�  ster ge�ffnet, mit dem Sie die Multimedia-datei abspielen k�   der Auswahl einer Multimedia-Datei wird dieses Kontrollfen�  EW.BMP /Macro /Play /Popup /Just L!�A/P /Just L /Text Nach�  /Just L!�R /I /Jump /Link E:\WORK\HINT_R~1.11\HELPFILE\MMVI�   �-�   !�' /T /Just L /Text Das Multimedia-Fenster!�
 /N �  n markiert. Wollen Sie einen Hinweis doch nicht lesen (viel    �                                                             ormalerweise das komplette Bild) angezeigt werden.  
� � �  er  �    �  	  � 4010   �  ��H�      � Fortschrit�  tsanzeige;Bilder;�� S�     � Das Bildanzeige Fenster���   b�     �  �� 	�5  o-�   !�( /T /Just L /Text Das Bil�  danzeige-Fenster!�
 /N /Just L!�S /I /Jump /Link E:\WORK\HI�  NT_R~1.11\HELPFILE\PICVIEW.BMP /Macro /Play /Popup /Just L!�  ter,(Global), 0,<Das Multimedia Fenster>!�3 neue Informatio�  �� /P /Just L /Text Die Anzeige unten rechts gibt den Forts�  chritt beim Laden des Bildes an. Mit Schlie�en verlassen Si�  e das Bildanzeige-Fenster. �ber die Auswahlliste k�nnen Sie     direkt zu verwandten Themen springen.  
� �             �  ie�en. �ber die Auswahlliste unten k�nnen Sie sofort zu ver�   k�nnen Sie das Fenster mit dem Close-Icon oben rechts schl�  leicht ist Ihnen ja inzwischen eine neue Idee gekommen), so    wandten Themen springen.  
� �                           �  n�s;�� E�     �	 Bedienung�� T�     �  �� 	��  -��     !�' /T /Just L /Text Hinweise zur Bedienung!�
 /N /Just�   L!�S /P /Just L /Text Wenn Sie The Hint Library starten, sQ  ehen Sie das folgende Fenster:!�6 /I /Link E:\WORK\HINT_R~1�  ?!�
 /N /Just L!�� /B /Just L /Text Neue Programmversionen,     �                                                        �  �  ��� 
� 0 7 P     � Topic@Lizenzvertrag  �  �    ���� 
v I P e   1  �, Topic@Eigenentwicklung von     >                                                         �  te festhalten und an die gew�nschte Position ziehen. 
.�  r Baumansicht bewegen, indem Sie sie mit der linken Maustas    ick �ffnen Sie das Informationsfenster.  
� �                ditors  
� �                                             �  �  ks�� 
� 9 @ Y   !  � Topic@Das Multimedia Fenste    uellen Thema hinzugef�gt.  
� �                          �    	  � 3000   �  ��:w   !  � Sprachen;Hauptfenster;Me�   werden!�b /B /Just L /Text Reader:��Mehrzeilige Darstell�  ung von Eintr�gen��Unterst�tzung f�r Verkn�pfungen!�� /B /J,  q  ���� 
� ) 0 I     � Topic@Inhalt  �    �  
  n,(Global), 0,<Das Infoedit Fenster>!�9 neuen Bildeintrag,(    INT LIBRARY !������  
� �                                �  mbers.aol.com/thlhome/index.htm����Viel Vergn�gen mit THE H�  ost.rwth-aachen.de����The Hint Library Homepage:��http://me�  l:   SMeier7777@aol.com oder��               Stefan.Meier@p�  , Erfstr. 65, 52249 Eschweiler��AOL:      SMeier7777��e-Mai�  rn o.�. erreichen Sie mich unter:��Post:       Stefan Meier�  ene THL-Dateien erstellen.����Bei Fragen, Anregungen, Fehle�   generiert.��Informationen hierzu finden Sie im Kapitel Eig�  t der "�bersetzer", der aus Ihren "Rohdaten" eine THL-Dateil  ust L /Text Editor:��Neues Editor-Design��Verschieben von�  �  ���� 
� , 3 L     � Topic@Bedienung  �    ��  arbeitet��Verkn�pfungen zwischen Eintr�gen k�nnen definiert�  ter werden die Informationen dargestellt (Nur-Lesen). Die A�  �  �r�� 
� 1 8 M     � Topic@Was ist neu...  �  �    �    �    �  ��?\     �  �� F�     � Was ist�   neu in Version 1.1�� U�     �  �� 	e�  �-�  
 !�- /T�   /Just L /Text Was ist neu in Version 1.1 ?!�
 /N /Just L!��  $ /H 1 /Just L /Text Entfernte Fehler:!�� /B /Just L /Text �  Allgemein:��Rechtschreibfehler in den Sprachpaketen korri�  giert��Ladefehler bei Bildern konnten Programmfehler verurs�  achen!�X /B /Just L /Text Reader:��Die Hinweiszeile im Re�  ader wurde z.T. nicht richtig gesetzt.!�� /B /Just L /Text �  Editor:��Manchmal wurden die Kn�pfe im Editor nicht richt�  ig gesetzt��Nachdem ein Eintrag nach unten bewegt wurde, wa�  r er nicht mehr selektiert!� /H 1 /Just L /Text Neu:!�� /B�   /Just L /Text Allgemein:��Neuer "Informations"-Typ f�r "�  Nicht"-Hinweis-Texte��THL-Format f�r mehr Flexibilit�t �ber   uswahlliste unten gibt Ihnen Zugriff auf verkn�pfte Themen.   geben Sie den Text Ihrer Information ein und einen optiona�  IT.BMP /Macro /Play /Popup /Just L!�� /P /Just L /Text Hier�  �  �o�� 
� < C \   $  � Topic@Die Bedienung des Edi�  tors  �    �  	  � 6000   �  ��J�   �  �� Schrifta�  rt;Autor;Titel;Themen;Bilder;Multimedia-Dateien;Hinweise;Fo�  rmate;Dateien bearbeiten;THL-Dateien;THR-Dateien;THL-Editor    �                                                          �  -  i�� 
� 6 = R     � Topic@Informationsfenster�    �    �  �� #    �  ��Da     �  �� K�     � Da�  s Informationsfenster�� Z�     �  �� 	j  w-�   !�( �  /T /Just L /Text Das Informationsfenster!�
 /N /Just L!�T /�  I /Jump /Link E:\WORK\HINT_R~1.11\HELPFILE\INFOVIEW.BMP /Ma�  cro /Play /Popup /Just L!�� /P /Just L /Text In diesem Fens     schlie�en.  
� �  � 6020                              �   Mit dem Schlie�en-Knopf rechts oben k�nnen Sie das Fenster"  len Titel. Wenn Sie keinen Titel angeben, erscheint sp�ter    eintragen;�� L�     � Verkn�pfungen definieren�� [�       �  �� 	��  �-�   !�) /T /Just L /Text Verkn�pfunge  n definieren!�
 /N /Just L!�S /I /Jump /Link E:\WORK\HINT_R  ~1.11\HELPFILE\LINKWND.BMP /Macro /Play /Popup /Just L!�a/  , 0,<Wo gibt es...>!�3 Verkn�pfungsfensters,(Global), 0,<Li  Das Themen Editierfenster, 0,!�- THL-Homepage nach,(Global)  l), 0,<Das Themen Editierfenster>!�3 Themen-Editierfenster,  obal), 0,<Das Hinweis Editierfenster>!�3 neues Thema,(Globa	  Global), 0,<Das Bilder Editierfenster>!�6 neuen Hinweis,(Gl  �  ��� 
� 7 > W     � Topic@Das Infoedit Fenster    �    �  	  � 6010   �  ��Ef     �  �� P�       � Das Infoedit Fenster�� _�     �  �� 	o�  P-�   !�  0 /T /Just L /Text Das Informations-Eingabefenster!�
 /N /J�  ust L!�T /I /Jump /Link E:\WORK\HINT_R~1.11\HELPFILE\INFOED    im Reader das Wort "Information".  
� �                     P /Just L /Text In diesem Fenster k�nnen sie zum aktuell in  �  ��� 
� < C \   $  � Topic@Das Bilder Editierfen^  ster  �    �  	  � 5010   �  ��J�   5  �0 Koordina     !�                                                            nks definieren>!�                                              seditor angezeigt.  
� �                                   kn�pfungen hinzuf�gen;Verkn�pfungen ver�ndern;Verkn�pfungen  rn definieren, wird immer der erste Eintrag aus dem Bereich  en Auswahllisten.��WICHTIG: Wenn Sie Verkn�pfungen zu Bilde   Solche Verkn�pfungen erscheinen dann sp�ter im Reader in d  . Mit dem "Zeile l�schen" - Knopf entfernen Sie eine Zeile.  ann eine Beschreibung f�r die Verkn�pfung eintragen sollten  . Es wird dann eine neue Zeile erzeugt werden, in der Sie d   den Zieleintrag aus der Baumansicht in dieses Fenster hier  ren. Um eine Verkn�pfung hinzuzuf�gen, "ziehen" Sie einfach   der Baumansicht selektierten Eintrag Verkn�pfungen definie"      �  	  � 6050   �  ��A�   \  �W Verkn�pfungen;Ver                                                               "                                                             #                                                             $                                                             %                                                             &                                                             '                                                             (                                                             )                                                             *                                                             +                                                             ,                                                             -                                                             .                                                             !    b��� 
� 3 : S     � Topic@Links definieren  �