���Z     @  W   I�      �   &                                       
    �                                                    !   �   ?s 	   ,          � Project@Options� -�   !�     7   \+ 	   -          � File@@Version2.1  � 1.1     (                                                          1   f   TOPIC VERSION OBJARRAY BROWSE_SEQUENCE BUILD_TAG CONTEX    link viewHandles 7                                            _ISECT_iterator _AE_Sorter _AE_mark _SysInfoFlags _outside_   Metafile VbPicture VbVarArray VeRec ViewEngine WinImage _AE   r VB_Historian VB_View VbCurrency VbDibBitmap VbFixArray Vb	   ng SystemDatabase TextFileDatabase TrashCollector TreeWalke
   Real RecordMark RuleSpecifier SchemaEngine SmartString Stri   adStream NamedData NamedMonad NilMonad Number Presentation    Dictionary Integer LogStream Monad MonadArray MonadFile Mon   tion Bcd36 Boolean ClassDesc ClassMethod ComboElement Date    Set AdRec AeAccessSet AgilityDatabase ArrayDatabase Associa   ]  YAccessCombo AccessEngine AccessItem AccessRule Accessh                   .       ,       )       8       	�     ..     E3     O�     P�     QI     S�     U�     W�     b�     k�     }�     ~�     ��     �r     ��     ��     �,     ��     ��     ��     ��     �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �0    !� BuildAll!� 0!� Inhalt!�$ � 1997 Stefan Meier, THL-Hi@   ump Der THL Reader /Link /Macro /Play /popup /Just L /Text "   ust L /Text General help on using The Hint Library!�Q /L /J�   192,192,192), 0!�3 "Index", ( 511, 0, 511, 1023), , , (192,$   , (192,192,192), 0!�4 "Glossary", ( 0, 0, 511, 1023), , , (%    511), , , (192,192,192), 0!�. "", ( 0, 511, 1023, 511), , &   4, 64, 832, 832), , , (192,192,192), 0!�, "", ( 0, 0, 1023,'   . "The Hint Library 1.1", , , , (192,192,192), 0!�- "", ( 6(   !  �� 	   -          � F1ProjectWindows�-�  t !�    �  !�  !�  !�  !�  !�                                      *     !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !+   �   �� 	   -          � F1ProjectButtonsZ -�   !�O  �C adding multimedia files,(Global), 0,<Das Multimedia Edit-   �    	   .          � F1ProjectGlossary�-�  # !     !� 0!� 0!� No!�  !� The Hint Library 1.1!� 1!�  !�  /   lfe 1.1.1!�  !�  !� E:\WORK\HINT_R~1.11\APP.ICO!� 0!�  !�"    T_STRING HELP_MACRO KEYWORDS TOPIC_TITLE NOTE              A    None , !�F Title , Arial ,  18 ,  120 ,  250 ,  40 ,  40 ,2   le , Arial ,  18 ,  120 ,  250 ,  40 ,  40 ,  0 , -1 ,  0 ,3   8 ,  120 ,  250 ,  40 ,  40 ,  0 , -1 ,  0 , None , !�F Tit4    ,  40 ,  40 ,  0 , -1 ,  0 , None , !�F Title , Arial ,  15    1 , -1 ,  0 , None , !�F Title , Arial ,  18 ,  120 ,  2506    Title , Times New Roman ,  24 ,  120 ,  250 ,  40 ,  40 , 7   @'  3 	 	  ,          � F1ProjectStyle2'-�  � !�P�   its!�P /L /Jump Lizenzvertrag /Link /Macro /Play /popup /Ju9   ump Referenzen /Link /Macro /Play /popup /Just L /Text Cred:   /Play /popup /Just L /Text What�s new in THL 1.1 ?!�C /L /J;   y /Popup /Just L /Text !�R /L /Jump Whats new /Link /Macro <    THL software and THL files ?!�1 /L /Jump /Link /Macro /Pla=   ... /Link /Macro /Play /popup /Just L /Text Where can I get>    /popup /Just L /Text The THL editor!�k /L /Jump Wo gibt es?   Reading THL files!�J /L /Jump Der Editor /Link /Macro /Play�P     0 , -1 ,  0 , None , !�R Paragraph , MS Sans Serif ,  10 Q   one , !�L Sub Heading , Arial ,  12 ,  180 ,  250 ,  40 ,  B    , Arial ,  12 ,  180 ,  250 ,  40 ,  20 ,  0 , -1 , -1 , NC    ,  250 ,  60 ,  20 ,  0 , -1 ,  0 , None , !�L Sub HeadingD   20 ,  0 , -1 ,  0 , None , !�H Heading , Arial ,  12 ,  180E    , None , !�H Heading , Arial ,  12 ,  180 ,  250 ,  60 ,  F   ding , Arial ,  12 ,  180 ,  250 ,  60 ,  20 ,  0 , -1 ,  0G   2 ,  180 ,  250 ,  60 ,  20 ,  0 , -1 ,  0 , None , !�H HeaH     60 ,  20 ,  5 , -1 ,  0 , None , !�H Heading , Arial ,  1I    None , !�R Heading , Times New Roman ,  24 ,  180 ,  250 ,J   ph , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 ,K    180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�J ParagraL     60 ,  0 ,  0 ,  0 , None , !�J Paragraph , Arial ,  10 , M    , None , !�J Paragraph , Arial ,  10 ,  180 ,  250 ,  20 ,N   raph , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0O   ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�J Parag`   20 ,  0 , -1 , -1 , None , !�L Sub Heading , Arial ,  12 , a    60 ,  0 ,  0 ,  0 , None , !�N Mono Spaced , Courier ,  10R   ne , !�N Mono Spaced , Courier ,  10 ,  180 ,  250 ,  20 , S   Courier ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , NoT    250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�N Mono Spaced , U     0 ,  0 , None , !�N Mono Spaced , Courier ,  10 ,  180 , V    Jump Label , Arial ,  10 ,  180 ,  250 ,  20 ,  20 ,  10 ,W     10 ,  180 ,  250 ,  20 ,  20 ,  10 ,  0 ,  0 , None , !�LX    20 ,  20 ,  10 ,  0 ,  0 , None , !�L Jump Label , Arial ,Y   ,  0 , None , !�L Jump Label , Arial ,  10 ,  180 ,  250 , Z   p Label , Arial ,  10 ,  180 ,  250 ,  20 ,  20 ,  10 ,  0 [    ,  180 ,  250 ,  20 ,  20 ,  10 ,  0 ,  0 , None , !�L Jum\    ,  20 ,  0 , -1 , -1 , None , !�L Jump Label , Arial ,  12]    , None , !�L Sub Heading , Arial ,  12 ,  180 ,  250 ,  40^   ding , Arial ,  12 ,  180 ,  250 ,  40 ,  20 ,  0 , -1 , -1_    180 ,  250 ,  40 ,  20 ,  0 , -1 , -1 , None , !�L Sub Heap    ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�N Monoq   10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�R Bib   60 ,  0 ,  0 ,  0 , None , !�Q Bitmap Paragraph , Arial ,  c    !�Q Bitmap Paragraph , Arial ,  10 ,  180 ,  250 ,  20 ,  d   ial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None ,e    20 ,  60 ,  0 ,  0 ,  0 , None , !�Q Bitmap Paragraph , Arf    None , !�Q Bitmap Paragraph , Arial ,  10 ,  180 ,  250 , g   ph , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 ,h    250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�Q Bitmap Paragrai   ,  0 ,  0 ,  0 , None , !�H Footnote , Arial ,  8 ,  180 , j   None , !�H Footnote , Arial ,  8 ,  180 ,  250 ,  20 ,  60 k   te , Arial ,  8 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , l     180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�H Footnom   0 ,  60 ,  0 ,  0 ,  0 , None , !�H Footnote , Arial ,  8 ,n    ,  0 , None , !�H Footnote , Arial ,  8 ,  180 ,  250 ,  2o    Spaced , Courier ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0�   tmap Jump Label , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  �   �R Enumerated Bullet , Arial ,  10 ,  180 ,  250 ,  20 ,  6r   l ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !s    ,  60 ,  0 ,  0 ,  0 , None , !�R Enumerated Bullet , Ariat    ,  0 , None , !�G Bullet , Arial ,  10 ,  180 ,  250 ,  20u   �G Bullet , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0v   l ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !w     250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�G Bullet , Ariax   60 ,  0 ,  0 ,  0 , Box , !�G Bullet , Arial ,  10 ,  180 ,y   0 , None , !�F Bullet , Arial ,  10 ,  180 ,  250 ,  20 ,  z   Label , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  {   ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�R Bitmap Jump |   0 ,  0 , None , !�R Bitmap Jump Label , Arial ,  10 ,  180 }   Jump Label , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  ~    180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�R Bitmap    0 ,  0 ,  0 , None , !�R Bitmap Jump Label , Arial ,  10 , �   0 ,  0 ,  0 ,  0 , None , !�R Enumerated Bullet , Arial ,  �    ,  10 ,  440 ,  250 ,  10 ,  10 ,  0 ,  0 ,  0 , None , !��     10 ,  10 ,  0 ,  0 ,  0 , None , !�M Outline Leaf , Arial�     0 , None , !�M Outline Leaf , Arial ,  10 ,  440 ,  250 ,�   ne Leaf , Arial ,  10 ,  440 ,  250 ,  10 ,  10 ,  0 ,  0 ,�   ,  180 ,  250 ,  10 ,  10 ,  0 ,  0 ,  0 , None , !�M Outli�   0 ,  0 ,  0 ,  0 , None , !�O Outline Branch , Arial ,  10 �   , !�O Outline Branch , Arial ,  10 ,  180 ,  250 ,  10 ,  1�   rial ,  10 ,  180 ,  250 ,  10 ,  10 ,  0 ,  0 ,  0 , None �    ,  10 ,  10 ,  0 ,  0 ,  0 , None , !�O Outline Branch , A�     0 , None , !�O Outline Branch , Arial ,  10 ,  180 ,  250�    Branch , Arial ,  10 ,  180 ,  250 ,  10 ,  10 ,  0 ,  0 ,�    180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�O Outline�   0 ,  0 ,  0 , None , !�R Enumerated Bullet , Arial ,  10 , �   umerated Bullet , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  �   10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�R En�   M Outline Leaf , Arial ,  10 ,  440 ,  250 ,  10 ,  10 ,  0�   tter Label , Arial ,  12 ,  180 ,  250 ,  20 ,  60 ,  0 , -�   180 ,  250 ,  20 ,  60 ,  0 , -1 ,  0 , None , !�S Index Le�   , -1 ,  0 , None , !�S Index Letter Label , Arial ,  12 ,  �    Letter Label , Arial ,  12 ,  180 ,  250 ,  20 ,  60 ,  0 �   ,  180 ,  250 ,  20 ,  60 ,  0 , -1 ,  0 , None , !�S Index�    0 , -1 ,  0 , None , !�S Index Letter Label , Arial ,  12 �   dex Letter Label , Arial ,  12 ,  180 ,  250 ,  20 ,  60 , �   10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�S In�   50 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�E Line , Arial ,  �    ,  0 ,  0 ,  0 , None , !�E Line , Arial ,  10 ,  180 ,  2�   0 , None , !�E Line , Arial ,  10 ,  180 ,  250 ,  20 ,  60�    Line , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  �   ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�E�     250 ,  10 ,  10 ,  0 ,  0 ,  0 , None , !�E Line , Arial �    ,  0 ,  0 , None , !�M Outline Leaf , Arial ,  10 ,  440 ,��   1 ,  0 , None , !�F Index , Arial ,  10 ,  180 ,  250 ,  20�    60 ,  0 ,  0 ,  0 , None , !�I Glossary , Arial ,  10 ,  1�    , None , !�I Glossary , Arial ,  10 ,  180 ,  250 ,  20 , �   abel , Arial ,  12 ,  180 ,  250 ,  20 ,  60 ,  0 , -1 ,  0�   0 ,  20 ,  60 ,  0 , -1 ,  0 , None , !�V Glossary Letter L�   None , !�V Glossary Letter Label , Arial ,  12 ,  180 ,  25�   l , Arial ,  12 ,  180 ,  250 ,  20 ,  60 ,  0 , -1 ,  0 , �     20 ,  60 ,  0 , -1 ,  0 , None , !�V Glossary Letter Labe�   e , !�V Glossary Letter Label , Arial ,  12 ,  180 ,  250 ,�    Arial ,  12 ,  180 ,  250 ,  20 ,  60 ,  0 , -1 ,  0 , Non�   0 ,  60 ,  0 ,  0 ,  0 , None , !�V Glossary Letter Label ,�    0 ,  0 , None , !�F Index , Arial ,  10 ,  180 ,  250 ,  2�   , !�F Index , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 , �   rial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None �   80 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�F Index , A�    ,  60 ,  0 ,  0 ,  0 , None , !�F Index , Arial ,  10 ,  1�   80 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�I Glossary �   ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�D Bar ,�    ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�D Bar , Arial ,  10 �   ,  0 ,  0 ,  0 , None , !�D Bar , Arial ,  10 ,  180 ,  250�   0 , None , !�D Bar , Arial ,  10 ,  180 ,  250 ,  20 ,  60 �   D Bar , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  �    ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !��     250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�F Image , Arial�   60 ,  0 ,  0 ,  0 , None , !�F Image , Arial ,  10 ,  180 ,�    0 , None , !�F Image , Arial ,  10 ,  180 ,  250 ,  20 ,  �    Image , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 , �   ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�F�    250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�F Image , Arial �     0 ,  0 ,  0 , None , !�I Glossary , Arial ,  10 ,  180 , �   ne , !�I Glossary , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,�   , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , Noj�    Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , Non�   ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,�   1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  �   e , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !��   !�;  , Arial ,  10 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 , Non�    ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , �   0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0�    0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  �   ,  0 ,  0 ,  0 , None , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 , �    ,  0 ,  0 , None , !�;  , Arial ,  10 ,  0 ,  0 ,  0 ,  0 �   ne , !�F Table , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0�   , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , No�     180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�F Table �    20 ,  60 ,  0 ,  0 ,  0 , None , !�F Table , Arial ,  10 ,�   ,  0 ,  0 , None , !�F Table , Arial ,  10 ,  180 ,  250 , �   e , !�F Table , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 "�     0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�;  , Arial ,  10 ,�    0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 , None , !�1  ,  ,  0 ,  0�    0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�;  , Arial ,  10 , �     0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 , �     ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,�    , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1�   �;  , Arial ,  10 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 , None�   ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�    ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 �   0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0�     0 ,  0 ,  0 , None , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  �     0 ,  0 ,  0 ,  , !�;  , Arial ,  10 ,  0 ,  0 ,  0 ,  0 ,�   ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,�    ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 �   0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0�     0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 , None , !�1  ,  ,  0 ,  ��    ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 �   e of the INIVISICLUES was to provide hints to several parts�   ch the idea of interactive providing hints. The main purpos�   ersions of the INVISICLUES(TM), but plane text does not mat�   inally the purpose of this software was to renew the INVISI�   CLUES(TM) in an electronical way to prevent the final loss �   of information. In addition there are different places in t�   he internet where you can find more or less complete text vm  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !� �   g /Link /Macro /Play /popup /Just L /Text Introduction and #   Overview!�a /L /Jump Bedienung /Link /Macro /Play /popup /J�   192,192), 0!�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  �  st L /Text Licence Agreement!�> /P /Just L /Text ������The      0 ,  0 ,  0 ,  , !�                                       �     0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 , �   ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,    of a game. These hints were divided into different topics   for further information.����Please remember: The sole inten�   ovide additional language support packs. Please contact me �   e help. I would be very pleased if anyone out there will pr�   ible shall be supported by the user interface and the onlin�    avaible to a wide range of users as many languages as poss�   s. (This is not limited to games !).��To make this software�   his project and develop their favourite hints to other user�    file collection. And everyone is invited to take part in t�   w the new purpose of The Hint Library is to build up a hint�   lso the capabilities to create new  hint collections. By no�   stem I decided not just to provide a read-only system but a�   elp as you need or as you wish. ����While developing the sy�   on with text-based solutions is that you just get as much h�   vided. The main advantage of these collections in comparisi�   while the hints were sorted due to the level of details pro�  t of this software is collecting information, It must not b  our raw data is invisible. ��Information about compiling yo  tion.��The compiler part, which generates a THL file from y  on on creating THL files please refer to The THL Editor sec  MP, JPEG, TARGA, PCX) in your files.��For further informati   text, multimedia files ( Sound, Videos ), and pictures ( B   collections with an easy to use interface. You can include   editor, which provides capabilites for creating new hint  se refer to Read THL-Files section.��The second part is the	  ia files( e.g. MIDI, AVI,...)��For further information plea
  the following types of hints: Text, pictures, and  multimed   receiving  of information shall be avoided. You will meet   t know explicitly requested information only. Inadvertandly  , provides capabilites for browsing hintfiles. You will ge  �Mainly there are two sections. The first one, ther Reader  e used for any commercial purposes.����About the software:�   u can find in Creating own THL files section.����Please sen  c/P /Just L /Text Author: Stefan Meier����Special thanks   :����Detlef Meister. Partially his MPICVIEW-Project is u  sed to display  PCX-,TGA- and JPEG-Files. Contact:��Meister  �  	  � 2000   �  ��;�   :  �5 Hint files;Infocom;Lang  uage files;Languages;Overview;�� F�     � Introduction  �� U�     �  �� 	��  �
-�   !�* /T /Just L /Text Intro�   duction and Overview!�
 /N /Just L!��
/P /Just L /Text Orig    .��  
� �                                                  ��The Hint Library 1.1 was created using Borland Delphi 2.0   made their adventures a milestone in computer history.����  @rz.fhtw-berlin.de����All former Infocom programmers, which  st L /Text The Hint Library 1.1!� /T /Just L /Text  Conten�   ts!�
 /N /Just L!� /P /Just L /Text !�U /L /Jump Einleitunw  an Meier, Erfstr. 65, 52249 Eschweiler��AOL:      SMeier777  d questions, announces or bug reports to:��Mail:       Stefj   	�M  �-�   !� /T /Just L /Text Credits!�
 /N /Just L!�#   of the notice.  Termination of the right to distribute doe$  s not affect distributors' other duties in this license.���%  �Many thanks go to Detlef Meister for his freeware project &  MPICVIEW. Parts of this project are used for displaying JPE'  G,TARGA and PCX files.��You can contact Detlef Meister at:�(  �Meister@rz.fhtw-berlin.de�� ��Enjoy The Hint Library!����C)  ontact:��Stefan Meier, Erfstr. 65, D-52249 Eschweiler, Germ*  any��AOL:��SMeier7777��E-Mail:��SMeier7777@aol.com��Stefan.    Meier@post.rwth-aachen.de��  
� �                        �  cture will be displayed. Ordinary the first hot spot contai  �  >;�� 
� - 4 M     � Topic@Einleitung  �    j  BMP /Macro /Play /Popup /Just L!�� /P /Just L /Text This wi/  V  i��� 
E - 4 I     � Topic@Referenzen  �    0  �    �    �  ��;�   1  �, Author;Borland Delphi;Greet!  ings;Information;�� B�     � Credits�� Q�     �  ��""   must stop distributing this archive 30 days after the date3  e to the ftp-Site given at the bottom of this document.����4  Distribution through retail and wholesale stores requires s5  pecific written permission.��Distribution through "magazine6  - compact disks" or "magazines-floppy disks" requires speci7  fic written permission.��No distributor may charge more tha8  n $8 US (or the appropriate value in other currencies, e.g.9   12 DM) for this archive.����Vendors' entire collection of :  THL files must be stored on a reasonably small number of di;  sks; distribution of hint files over excessive numbers of d<  isks is prohibited.  No more than $8 US (or the appropriate=   value in other currencies, e.g. 12 DM) may be charged for >  any disk containing THL files.��These terms are a condition?   of distribution of this archive and apply to all THL files@   written by any hint author.����Right to distribute this ar1  chive may be terminated by written notice, and distributors�2  ase send a copy to me. The easiest way is to upload the filC   documentation are provided "AS IS" and without warranty ofD   any kind and the author expressly disclaims all other warrE  anties,��express or implied, including, but not limited to,F   the implied warranties of merchantability and fitness for G  a particular purpose. Under no circumstances shall Stefan MH  eier be liable for any incidental, special or consequentialI   damages that result from the use or inability to use the sJ  oftware or related documentation, even if Stefan Meier has K  been advised of the possibility of such damages.����If you L  intent to write THL-files with the included editor and distM  ribute them you should always contact me to tell me about yN  our project and check out if anyone else is working on a hiO  nt file for the given game. Although the use of the softwarP  e is free you are NOT ALLOWED to take charge for your indivA  idual THL-files.  If you want to spread your THL-Files, ple�B  is software in your possession.����The software and relatedS  ement between you and Stefan Meier covering your use of TheT   Hint Library. Be sure to read the following agreement befoU  re using the software. IF YOU DO NOT AGREE TO THE TERMS OF V  THIS AGREEMENT, DO NOT USE THE SOFTWARE AND DESTROY ALL COPW  IES OF IT.��This copyright software is distributed as freewX  are. You may use this software without any charge and may dY  istribute to others. The software is owned by Stefan Meier Z  and is protected by FR Germany copyright laws and internati[  onal treaty provisions. Therefore, you must treat the softw\  are like any other copyrighted material (e.g., a book or mu]  sical recording).����You may not rent or lease the software^  , nor may you modify, adapt, translate, reverse engineer, d_  ecompile, or disassemble the software.��If you violate any `  part of this agreement, your right to use this software terQ  minates automatically and you then destroy all copies of thR  ment!�
 /N /Just L!�(/P /Just L /Text This is a legal agrec   exists The Hint Library��!�{ /R /Link E:\WORK\HINT_R~1.11\d  HELPFILE.GB\EDITOR~1.BMP /Just L /Text Editor opens the ee  ditor window with a blank formular.!��/R /Link E:\WORK\HINf  T_R~1.11\HELPFILE.GB\SPRACH~1.BMP /Just L /Text Use Languag  ge - Select language to open a dialog for choosing a languh  age support package. By default only the English language pi  ackage is included, but the system can easily be extended. j  For additional language packages please refer to THL homepak  ge. WithLanguage - Save language setting you can decide i�  f the chosen language will be selected each time you start �  files;Title;Topics;�� U     � Using the THL editor�� �   !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�o    �  	  � 7000   �  ��>�   +  �& Conditions;License;Dp  istribution rules;�� I�     � Licence Ageement�� X�  a     �  �� 	�&  f-�   !�" /T /Just L /Text Licence Agree�b  oosing a THL file by title and opening the Reader..��Exits  xt Open a THL file for reading hints. Information on readint  g hints you cam find in the THL Reader section.!�� /R /Linku   E:\WORK\HINT_R~1.11\HELPFILE.GB\VOPEN.BMP /Just L /Text Opv  en a THL file in verbose mode. You will not see the filenamw  es but the titles of the THL files.!�U /R /Link E:\WORK\HINx  T_R~1.11\HELPFILE.GB\EXISTF~1.BMP /Just L /Text Opens the ey  ditor.!�T /R /Link E:\WORK\HINT_R~1.11\HELPFILE.GB\HELP.BMPz   /Just L /Text Open this help file.!�� /R /Link E:\WORK\HIN{  T_R~1.11\HELPFILE.GB\INFO.BMP /Just L /Text Show program in|  formation like program version and contact information.!�U }  /R /Link E:\WORK\HINT_R~1.11\HELPFILE.GB\EXIT.BMP /Just L /~  Text Exit The Hint Library!�& /H 2 /Just L /Text The progra  m menues:!�� /R /Link E:\WORK\HINT_R~1.11\HELPFILE.GB\DATEI�  M~1.BMP /Just L /Text Select File open for choosing a THLq   file and opening the Reader.��Select Verbose open for ch"r  ink E:\WORK\HINT_R~1.11\HELPFILE.GB\OPENBTN.BMP /Just L /Te�    	  � 3000   �  ��:x   "  � Main window;Menues;Langu�  gram version, contact adresses and other usefull informatio�   brings up an information dialog where you can find the pro�  s you instructions on using the Windows help system��Info�  search the helpfiles by key words��Help - Using help show�  nline help and go to contents page��Use Help - Search to �  HILFEM~1.BMP /Just L /Text Use Help - Contents to start o�  automatically.!��/R /Link E:\WORK\HINT_R~1.11\HELPFILE.GB\�  ages;�� E�     � Operating instructions�� T�     �  �  �� 	��	  �-�   !�' /T /Just L /Text Operating instructio�  ns!�
 /N /Just L!�Y /P /Just L /Text After starting The Hin�  t Library you will encounter the following window:!�9 /I /L�  ink E:\WORK\HINT_R~1.11\HELPFILE.GB\MAIN.BMP /Just L!� /H     Hint Library � 1996-97 Stefan Meier  
� �                �  /Just L /Text !�  /H 2 /Just L /Text Speedbuttons:!�� /R /L"�  �	  ���� 
} , 3 L     � Topic@Bedienung  �    �l  t;Hints;Multimedia files;Pictures;THL Editor;THL files;THR �  inks;informations;Author;Edit files;Editor;File formats;Fon�  tors  �    �  	  � 6000   �  ��J�   �  �� Define l�  {  ���� 
� < C \   $  � Topic@Die Bedienung des Edi�  L!�r /L /Jump Was sind THL Dateien... /Link /Macro /Play /p�    �-�   !� /T /Just L /Text The THL editor!�
 /N /Just �  iles,edit;�� F�     �
 The editor�� U�     �  �� 	�H�  �  	  � 5000   �  ��;}   &  �! Editor;THL Editor;THL f�  N  8��� 
� ) 0 I     � Topic@Inhalt  �    �  �  _  s�� 
U : A Z   "  � Topic@Das Bildanzeige Fenst�    �  	  � 4000   �  ��?}   "  � Read hints;Reader;T�  HL Reader;�� J�     � The THL Reader�� Y�     �  ���  x  ��� 
P 9 @ Y   !  � Topic@Das Multimedia Fenste-  !�V /I /Jump /Link E:\WORK\HINT_R~1.11\HELPFILE.GB\INFOWND.    e hint file.  
� �                                            recommened due to compability reasons.  
� �            �  t L /Text Eventually save your data as THR-File (highly rec�  ommened). A THR-File saves your data without compiling them�  .��CAUTION: THL-File can not be edited with the THL-Edito�  r anymore. Always keep a copy of your THR-File at a save pl�  ace.!�9 /B /Just L /Text Compile the editor data into a THL�  -File.!� /H 1 /Just L /Text !�2 /H 1 /Just L /Text The str�  ucture of THR/THL-Files:!�� /P /Just L /Text Ordinary a hin�  t collection is divided into deveral topics. These topic co�  ntain subtopics or hints.There are different hint types:!�2�   /B /Just L /Text Text ( single or multiple lines )!�� /B /�  Just L /Text Pictures, supported file formats: Bitmap, JPeg�  , PCX, Targa��Special features: You may define parts of pic�  tures and attach independent descriptions.!�� /B /Just L /T�  ext Multimedia-Files, suported formats: WAV, AVI, MIDI, MOV�  . Some additional formats are supported, but the use is not��  hints, include pictures, ... with the THL-Editor!�� /B /Jus�  opup /Just L /Text What are THL files, how are they created^  ster  �    �  	  � 5010   �  ��J�   3  �. Areas;Co�  C  w��� 
� 3 : S     � Topic@Links definieren  ��      �  	  � 6050   �  ��A�   2  �- Links;Adding link�  s;Defining links;Edit links;�� L�     � Defining links�  *  J�� 
� : A V   "  � Topic@Was sind THL Dateien.�  ..  �    �    �    �  ��H�   F  �A Pictures;File �  formats;Hints;Multimedia files;THL files;THR files;�� O� �      � What�s a THL-File ?�� ^�     �  �� 	�!  =-�  �   !� /T /Just L /Text THL-Files!�
 /N /Just L!�/P /Just �  L /Text THL-Files are binary files which contain text, pict�  ures and multimediadata. They are designed for the use with�   the "reader" of this software, but they are not suitable f�  or ordinary texteditors. In general the creation of THL-Fil�  es consists of three main steps:!�G /B /Just L /Text Enter �  ?!�u /L /Jump Eigenentwicklung von Hinweissammlungen /Link �  the progress of the THL project.!�� /B /Just L /Text Think �   one topic and to make it possible to me to keep an eye on �  ile about your topic. This is done to avoid double works on�  should contact me to check if anyone else is working on a f�  advices:!� /B /Just L /Text Before starting your work you �  wn hint collections, please pay attention to the following �  st L!�v /P /Just L /Text If you wish to design and spread o�   !�, /T /Just L /Text Creating your own THL files!�
 /N /Ju�   Userdefined files;Development;THL files;�� ^�   !  � Cr�  Hinweissammlungen  �    �    �    �  ��W�   -  �(�  �  �j�� 
. I P e   1  �, Topic@Eigenentwicklung von �  eation of hint collections�� m�     �  �� 	��  �-�  	�  Q  �:�� 
b - 4 M     � Topic@Der Editor  �    4  les.!�l /L /Jump Die Bedienung des Editors /Link /Macro /Pl�  /Macro /Play /popup /Just L /Text Development of own THL fij�  about the structure of your hint collection. Where can ques�  ernativly you can send the file by mail or name a internet �  ng ftp-site:��ftp://members.aol.com/thlhome/incoming��Alt�   The easiest way to do is uploading the file to the followi�  /B /Just L /Text Please send a copy of your THL file to me.�  lace. A THL file can not be edited with the THL editor.!��  file, but always keep a copy of your THR file at a secure p�  ly. Remember that anyone is able to edit the data in a THR �  riginal.!�� /B /Just L /Text You should spread THL files on�  doubt about legimitation please contact the author of the o�  mmercial hint books into electronical systems. If you have �  any copyrights. Ordinarily it is prohibited to transform co�  sions.!�� /B /Just L /Text Please make sure not to violate �  solution with different solutions to prevent errors or omis�  al parts can be defined ?!�_ /B /Just L /Text Compare your �  tions occur ? When is picture support usefull ? Which logic�    site where I can download the file.  
� �                �   I get...?�� X�     �  �� 	�{  �-�   !�% /T /Just L �  /Text Where can I get... ?!�
 /N /Just L!�| /B /Just L /Tex�  t New program versions, language support packages, and THL �  files:��http://members.aol.com/thlhome/index.htm!�� /B /J�  ust L /Text If you prefer FTP try this:����THL software:���  a  U��� 
~ 1 8 Q     � Topic@Der THL Reader  �  `    !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !     � Contents�� Q�     �  �� 	sE  �-�   !�% /H /Ju�  Reader,(Global), 0,<Der THL Reader>!�- THL-Homepage nach,(G�  Themen-Editierfenster,Das Themen Editierfenster, 0,!�' THL n  /  6�� 
� 0 7 P     � Topic@Lizenzvertrag  �  �  ext Bugs removed:!�g /B /Just L /Text General:��Spelling �  errors corrected ��Load errors on pictures caused malefunct�  ions��!�V /B /Just L /Text Reader:��The hint line of the �  reader window was not set correctly��!�� /B /Just L /Text "�  ks;New program versions;THL files;�� I�     � Where can    ft mouse button pressed. 
)9                          1   /P /Just L /Text PLEASE PAY ATTENTION TO THE ADVICES ON CR�  ~1.11\HELPFILE.GB\EDITOR.BMP /Macro /Play /Popup /Just L!�L�  e THL editor!�
 /N /Just L!�U /I /Jump /Link E:\WORK\HINT_R�  e info edit window>!�9 new picture links,(Global), 0,<Das B�  to delete the currently selected line.��IMPORTANT: If you d�  Text What�s new in THL 1.1!�
 /N /Just L!�  /H 1 /Just L /T�  ilder Editierfenster>!�1 new topic,(Global), 0,<Das Themen �  Editierfenster>!�< picture display window,(Global), 0,<Das ?  ultimedia Fenster>!�; Multimedia-Editierfenster,Das Multime    n.  
� �                                                 k  s:��ftp://members.aol.com/smeier7777/thl_lang����THL file�  ftp://members.aol.com/nicetoon/thl1.gb����Language package�  	  � 1000   �  ��7j     � Contents;Overview;�� B�      !�  !�                                                     "�  em and move it to the desired location while keeping the le  Reader to display the title of your document. Please note t  hat the use non standard fonts may cause unwanted  effects   on computer system which do not have the fonts installed.!�  � /E /Just L /Text Use this window to enter copyright notic  e, e.g. Written 1997 by Harry Hummel. This field must be   filled in for proper compilation.!�N /E /Just L /Text Here 	  you can enter additional information about your project.!�
   /P /Just L /Text !� /H 1 /Just L /Text The menues:!�� /P   /Just L /Text Use the File - menu to save your project as   THR-File and to close the editor.��Use the Project -menu   to compile your work into the THL format!�- /H 1 /Just L /  Text Additional functionallity:!�/P /Just L /Text Clickin  g the right mouse button in the tree view opens a popup men  u for faster access to creation functions.��You can move en  tries within the tree view with drap and drop. Select an it  s button you can choose a font which will be used with the   w information to your project.!�� /E /Just L /Text This but  ton opens the link editor where you can define references t  o related entries in your file.��Refer to Links section for   instructions.!�� /E /Just L /Text Edit the selected entry.   The software will select the appropriate window for the en  try. It is not possible to change type of an entry.!�� /E /  Just L /Text This buttons moves the currently selected item   within its level upwards. Associated children will be move  d either.!�$ /E /Just L /Text Moving downwards...!�� /E /Ju  st L /Text Delete the currently selected entry. Please note   that you even delete all children of this entry. Use this   function carefully !!�� /E /Just L /Text Enter a title for   your document here. This is not a file name, but a title wh   ich appears as header in the Reader. This entry is nessesar  y for successfull compilation.!�/E /Just L /Text With thi�  ifferent systems.!�D /E /Just L /Text Here you can add a ne#   your current project. Hints are marked with the prefix HIN$  T, pictures are marked with PIC, information is marked with%   INFO, and multimedia files are marked with MM. You always &  will see the starting characters of a title.!�[ /E /Just L '  /Text Pressing this button open a window for adding a new t(  opic to your project.!�� /E /Just L /Text This button opens)   the picture editor which is used to add new picture links *  or area definitions to your project.!�= /E /Just L /Text He+  re you can add a new hint to your project.!��/E /Just L /T,  ext Pressing button no 5 open a window for adding multimedi-  a files to your project. Please note that normally video fi.  les are rather large and therefore the size of the THL file/   will increase significantly. Although the multimedia suppo0  rt of THE HINT LIBRARY only depends on the capabilites of y!  our system, unusual files formats may not be supported by d�"  EATING THL FILES !!�/E /Just L /Text This tree view showsA  ster  �    �  	  � 5030   �  ��J~     � Text;Add2  �  )j�� 
O < C \   $  � Topic@Das Themen Editierfen�  ay /popup /Just L /Text Instructions on using the editor. 6  pe for non-hint-information��Restructured file format for m7  ore flexibility��Direct links between entries can be defini;  ed��!�L /B /Just L /Text Reader:��Multiple line support��    e��  
� �                                                8  nhanced Save/Compile - Menu��Save file check on editor clos9  w editor design��Moving editor entries via drag and drop��E:  Added support for links��!�� /B /Just L /Text Editor:��Ne�   Reader>!�# Reader,(Global), 0,<Der THL Reader>!� Reader:,�   Hinweis Editierfenster>!�2 new information,(Global), 0,<Th=  l), 0,<Das Multimedia Fenster>!�1 new hint,(Global), 0,<Das>  dia Editierfenster, 0,!�? Multimedia-Kontrollfenster,(Globa�  r  �    �  	  � 6020   �  ��Gh     �  �� R�   P  ing topics;�� U�     � The topic edit window�� d�   �  u close the window with the OK button the new hint will be B  /P /Just L /Text Enter your text into the Text field. If yoC  11\HELPFILE.GB\HINTEDIT.BMP /Macro /Play /Popup /Just L!�� D  it window!�
 /N /Just L!�W /I /Jump /Link E:\WORK\HINT_R~1.E       �  �� 	��  (-�   !�% /T /Just L /Text The hint edF  ding hints;Text;�� V�     � The hint edit window�� e�G  nster  �    �  	  � 5020   �  ��K�     � Hint;AdH  �  mM�� 
S = D ]   %  �  Topic@Das Hinweis Editierfe    c will be added to your project.  
� �                   J  . If you close this window with the OK button, the new topiK  Just L /Text Enter the title of your topic at the TEXT lineL  HELPFILE.GB\TOPEDIT.BMP /Macro /Play /Popup /Just L!�� /P /M  window!�
 /N /Just L!�V /I /Jump /Link E:\WORK\HINT_R~1.11\_  ierfenster>!�: Bild-Anzeigefenster.,(Global), 0,<Das BildanN    �  �� 	��  6-�   !�& /T /Just L /Text The topic edit �  is-Anzeigefenster,(Global), 0,<Das Hinweis Fenster>!�* Hinwa  hould edit the description or remove the item.��If you closR  ure will be added to the hotspot list automatically. Show sS  a description. On selecting a new picture the complete pictT  l be added to the hotspot list. Now you just have to enter U  use. On releasing the left mouse button the marked area wilV  ton into the picture and marked the area by dragging the moW  e separate picture areas: Click and hold the left mouse butX  filename at the FILE field. Use the hotspot editor to definY  ro /Play /Popup /Just L!�-/P /Just L /Text Please enter a Z  Jump /Link E:\WORK\HINT_R~1.11\HELPFILE.GB\PICEDIT.BMP /Mac[  /Just L /Text The picture edit window!�
 /N /Just L!�V /I /\  icture edit window�� d�     �  �� 	��  �-�   !�( /T ]  ordinates;Pictures;Progress indicator;�� U�     � The ph  zeige Fenster>!�1 Bild-Editierfenster,Das Bilder Editierfen�  �  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  p  e the window with the OK button, the new entry will be addeq  /Play /Popup /Just L!�� /P /Just L /Text Please enter a filb  mp /Link E:\WORK\HINT_R~1.11\HELPFILE.GB\MMEDIT.BMP /Macro c   L /Text The multimedia edit window!�
 /N /Just L!�U /I /Jud  a edit window�� h�     �  �� 	�u  �-�   !�+ /T /Juste   description;Multimedia files;�� Y�     � The multimedif  rfenster  �    �  	  � 5040   �  ��N�   '  �" File}  ster, 0,!�S Creating own THL files section,(Global), 0,<Eig�  wn list provides access to related topics. Use upper right i  ndow displays the information text (read-only). The drop do    s:��ftp://members.aol.com/smeier7777/thlfiles��  
� �      be displayed.   
� �                                     l  e links to this picture always the first hotspot area will m  eparate entries for the THL files.��IMPORTANT: If you definn  y per picture in your project, the compiler will generate so  d to your project. Although you only will see a single entr"�  ename in the File field or choose a file with the Browse bus  .  �(�� 
� , 3 H     � Topic@Whats new  �    ��      �    �  ��:W     �  �� A|     � What�s new i    /thlhome/index.htm����Enjoy THE HINT LIBRARY !��  
� �   t  ftp://members.aol.com/thlhome��oder��http://members.aol.comu  n.Meier@post.rwth-aachen.de����The Hint Library Homepage:��v  7��e-Mail:   SMeier7777@aol.com oder��                Stefa�  �' Der-THL-Editor,(Global), 0,<Der Editor>!� editor,(Globax  weissammlungen>!�' Der THL-Editor,(Global), 0,<Der Editor>!5  tures:!�� /B /Just L /Text General:��Added information tyy  ating your own files.,(Global), 0,<Eigenentwicklung von Hin{  (Global), 0,<Eigenentwicklung von Hinweissammlungen>!�M Cre|  enentwicklung von Hinweissammlungen>!�G CREATING THL FILES,     button adds the new entry to your project.  
� �        ~  t at the descriptiion field. Closing the window with the OK  tton. Afterwards enter a description f�r the multimedia hin��  \HELPFILE.GB\INFOEDIT.BMP /Macro /Play /Popup /Just L!�� /P�  e file. Double-clicking an item opens the specific topic. T�  here will will either encounter different subtopics or hint�  s:!�� /R /Link E:\WORK\HINT_R~1.11\HELPFILE.GB\HINTPIC.BMP �  /Just L /Text Text hints: Double-clicking a hint item opens�   the hint window. Because hints are sorted to their level o�  f detail a warning will raise if you try to read hint no 3 �  before hint no 2.!�� /R /Link E:\WORK\HINT_R~1.11\HELPFILE.�  GB\MMPIC.BMP /Just L /Text Multimedia hints: Double-clickin�  g a multimedia item brings up a multimedia control panel..!�  �� /R /Link E:\WORK\HINT_R~1.11\HELPFILE.GB\PICPIC.BMP /Jus�  t L /Text Picture hints: Double-clicking a picture item ope�  ns the picture display window.!�� /R /Link E:\WORK\HINT_R~1�  .11\HELPFILE.GB\INFOPIC.BMP /Just L /Text Information text:�   Double-clicking an information item opens the information     display window.  
� �                                    ��  tred in the window displays the main topics contained in th�    � The multimedia control panel�� a�     �  �� 	�o  �  edia files;Multimedia contral;Multimedia player;�� R�   !�  l), 0,<Der Editor>!�/ Editor:,(Global), 0,<Die Bedienung de�   pressing the Close icon in the upper right corner. The dro�  p down list provides direct access to related entries of th    e hint file.  
� �                                       �   !�' /T /Just L /Text The information window!�
 /N /Just L@  �  ���� 
� 9 @ Y   !  � Topic@Das_Infoanzeigefenste�  �  c�� 
k 0 7 P     � Topic@Wo gibt es...  �  �  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !� �   	�X  �-�  	 !� /T /Just L /Text The THL Reader!�
 /N /J�  ust L!�e /P /Just L /Text After opening and compilation of �  a THL file you will encounter the following window:!�U /I /�  Jump /Link E:\WORK\HINT_R~1.11\HELPFILE.GB\READER.BMP /Macr�  o /Play /Popup /Just L!�� /P /Just L /Text The list box cen��  �-�   !�- /T /Just L /Text The multimedia control panel!��  TVIEW.BMP /Macro /Play /Popup /Just L!��/P /Just L /Text A�  fter selecting a hint you will encounter the following wind�  ow. For reading the hint you have to click the SHOW HINT bu�  tton. After reading the hint you can close the window by pr�  esing the close button. This hint will be marked as "read".�   ��If you decide not to read the hint yet, you can abort by�  enentwicklung von Hinweissammlungen>!�N ERSTELLEN VON THL-D�  s Editors>!�Q Eigene THL-Dateien erstellen,(Global), 0,<Eig�    � The information window�� a�     �  �� 	q�  K-�      ides direct access to related topics.  
� �              �  nd stops a currently running media. The drop down list prov�   panel is shown. Pressing the OK button closes the window a�  ext After selecting a multimedia hint the following control�  .GB\MMVIEW.BMP /Macro /Play /Popup /Just L!�� /P /Just L /T�  
 /N /Just L!�U /I /Jump /Link E:\WORK\HINT_R~1.11\HELPFILE�  ust L!�W /I /Jump /Link E:\WORK\HINT_R~1.11\HELPFILE.GB\HIN    added to your project.  
� �                                 close button to hide the window.  
� �                   �  drop down list offers direct access to related topics in th�  . Pressing the Close button exists the display window. The �   lower left corner shows refers to the file loading process�  p /Just L!�� /P /Just L /Text The progress indicator in the�  WORK\HINT_R~1.11\HELPFILE.GB\PICVIEW.BMP /Macro /Play /Popu�  ATEIEN,(Global), 0,<Eigenentwicklung von Hinweissammlungen>�   picture display window!�
 /N /Just L!�V /I /Jump /Link E:\�  w�� b�     �  �� 	�V  �-�   !�+ /T /Just L /Text The�  rogress indicator;�� S�     � The picture display windo�  er  �    �  	  � 4010   �  ��H�   !  � Pictures;P�    �    �  	  � 4020   �  ��D{     � Hidden hint;Sh�  ow hint;�� O�     � The hint window�� ^�     �  �� �  	�  R-�   !�  /T /Just L /Text The hint window!�
 /N /J�    �"�� 
W 6 = V     � Topic@Das Hinweis Fenster�  ,(Global), 0,<Links definieren>!�$ Links,(Global), 0,<Links�   window,(Global), 0,<Das_Infoanzeigefenster>!�* link editor�  nster,Das Hinweis Editierfenster, 0,!�? information display�  eis-Dateien-lesen,(Global), 0,<(None)>!�5 Hinweis-Editierfe+  efine links to a picture, the first hot spot area of the pi�  �  `��� 
� < C \   $  � Topic@Das Bilder Editierfen�  d0    �  �� 	r  7-�   !�% /T /Just L /Text Using th�  n THL 1.1�� P�     �  �� 	`%  �-�  
 !�& /T /Just L /�  Editor:��Sometimes button states in the editor window are �  not set correctly��After moving down an entry in the editorz   the entry was not selected��!�  /H 1 /Just L /Text New fea<  Bildanzeige Fenster>!�+ Read THL-Files,(Global), 0,<Der THL     
� �                                                     �  r  �    �  	  � 4030   �  ��G�   @  �; Play multimg  ~  =%�� 
Q @ G `   (  �# Topic@Das Multimedia Editie�   definieren>!�= multimedia control panel,(Global), 0,<Das M�  l contain a "This is a sample link" entry whenever you sele�  ct the "This is a topic" topic. Use the delete line button �    �  	  � 8000   �  ��>�   ;  �6 Language support pacQ  !�. hint window.,(Global), 0,<Das Hinweis Fenster>!�8 Hinwe�  (Global), 0,!�' The THL editor,(Global), 0,<Der Editor>!�3 �  �  ��� 
� 7 > W     � Topic@The info edit window�    �    �  	  � 6010   �  ��Ez     � information e�  diting;�� P�      � The information edit window�� _�  �     �  �� 	��  0-�   !�% /T /Just L /Text The info edit�   window!�
 /N /Just L!�W /I /Jump /Link E:\WORK\HINT_R~1.11    er will state "information".  
� �                       �  ry. The title is optional. If no title is provided the read�   /Just L /Text Use this window to create an information ent    ns the complete picture.  
� �                           �   !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !���  In this example the drop down list of the reader window wil                                                               �                                                             �                                                             �                                                                 lobal), 0,<Wo gibt es...>!�                                      !�  !�  !�  !�  !�  !�  !�  !�  !�                       �  �� [�     �  �� 	�:  r-�   !� /T /Just L /Text Defin�  ing links!�
 /N /Just L!�V /I /Jump /Link E:\WORK\HINT_R~1.�  11\HELPFILE.GB\LINKWND.BMP /Macro /Play /Popup /Just L!��/�  P /Just L /Text This window displays all links definied for�   an entry. To add a new link, please mark the related entry�   in the tree view, and drag and drop it to this window. A n�  ew line will be added and you can enter a description for t�  he link. Later in the reader these links will apear in the �  associated drop down lists whenever the owner is selected. 