���Z     @  E   I�      �   &                                       
                                                        !   �   �6 	   ,          � Project@Options� -�   !�     7   \+ 	   -          � File@@Version2.1  � 1.1     (                                                          1   f   TOPIC VERSION OBJARRAY BROWSE_SEQUENCE BUILD_TAG CONTEX    link viewHandles 7                                            _ISECT_iterator _AE_Sorter _AE_mark _SysInfoFlags _outside_   Metafile VbPicture VbVarArray VeRec ViewEngine WinImage _AE   r VB_Historian VB_View VbCurrency VbDibBitmap VbFixArray Vb	   ng SystemDatabase TextFileDatabase TrashCollector TreeWalke
   Real RecordMark RuleSpecifier SchemaEngine SmartString Stri   adStream NamedData NamedMonad NilMonad Number Presentation    Dictionary Integer LogStream Monad MonadArray MonadFile Mon   tion Bcd36 Boolean ClassDesc ClassMethod ComboElement Date    Set AdRec AeAccessSet AgilityDatabase ArrayDatabase Associa   ]  YAccessCombo AccessEngine AccessItem AccessRule Accessh �                   .       ,       )       8       	�     ��     ��     �^     ��     ��     �~     ��     �J     ��     	�     
�     1     ,     �     -     �     �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           �0    !� BuildAll!� 0!� Inhalt!�$ � 1996 Stefan Meier, THL-Hi#    /popup /Just L /Text The THL editor!�k /L /Jump Wo gibt es�   ... /Link /Macro /Play /popup /Just L /Text Where can I get�   192,192,192), 0!�3 "Index", ( 511, 0, 511, 1023), , , (192,$   , (192,192,192), 0!�4 "Glossary", ( 0, 0, 511, 1023), , , (%    511), , , (192,192,192), 0!�. "", ( 0, 511, 1023, 511), , &   4, 64, 832, 832), , , (192,192,192), 0!�, "", ( 0, 0, 1023,'   . "The Hint Library 1.0", , , , (192,192,192), 0!�- "", ( 6(   �  *Q 	   -          � F1ProjectWindows�-�  Y !�    �  !�  !�  !�  !�  !�                                      *     !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !+   �   �� 	   -          � F1ProjectButtonsZ -�   !�O  �: Bild-Anzeigefenster.,(Global), 0,<Das Bildanzeige Fenste-   �  dx 	   .          � F1ProjectGlossary~-�   !   � 0!� 0!� No!�  !� The Hint Library 1.0!� 1!�  !�  !� /   lfe 1.0.1!�  !�  !� E:\WORK\HINT_R~1\APP.ICO!� 0!�  !�  !"    T_STRING HELP_MACRO KEYWORDS TOPIC_TITLE NOTE              A    None , !�F Title , Arial ,  18 ,  120 ,  250 ,  40 ,  40 ,2   le , Arial ,  18 ,  120 ,  250 ,  40 ,  40 ,  0 , -1 ,  0 ,3   8 ,  120 ,  250 ,  40 ,  40 ,  0 , -1 ,  0 , None , !�F Tit4    ,  40 ,  40 ,  0 , -1 ,  0 , None , !�F Title , Arial ,  15    1 , -1 ,  0 , None , !�F Title , Arial ,  18 ,  120 ,  2506    Title , Times New Roman ,  24 ,  120 ,  250 ,  40 ,  40 , 7   @'  3 	 	  ,          � F1ProjectStyle2'-�  � !�P:      � Contents�� Q�     �  �� 	s�  O-�   !�% /H /Ju;   st L /Text The Hint Library 1.0!� /T /Just L /Text  Conten<   ts!�
 /N /Just L!� /P /Just L /Text !�U /L /Jump Einleitun=   g /Link /Macro /Play /popup /Just L /Text Introduction and >   Overview!�a /L /Jump Bedienung /Link /Macro /Play /popup /J?   ust L /Text General help on using The Hint Library!�Q /L /J@   ump Der THL Reader /Link /Macro /Play /popup /Just L /Text "   Reading THL files!�J /L /Jump Der Editor /Link /Macro /Play�P     0 , -1 ,  0 , None , !�R Paragraph , MS Sans Serif ,  10 Q   one , !�L Sub Heading , Arial ,  12 ,  180 ,  250 ,  40 ,  B    , Arial ,  12 ,  180 ,  250 ,  40 ,  20 ,  0 , -1 , -1 , NC    ,  250 ,  60 ,  20 ,  0 , -1 ,  0 , None , !�L Sub HeadingD   20 ,  0 , -1 ,  0 , None , !�H Heading , Arial ,  12 ,  180E    , None , !�H Heading , Arial ,  12 ,  180 ,  250 ,  60 ,  F   ding , Arial ,  12 ,  180 ,  250 ,  60 ,  20 ,  0 , -1 ,  0G   2 ,  180 ,  250 ,  60 ,  20 ,  0 , -1 ,  0 , None , !�H HeaH     60 ,  20 ,  5 , -1 ,  0 , None , !�H Heading , Arial ,  1I    None , !�R Heading , Times New Roman ,  24 ,  180 ,  250 ,J   ph , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 ,K    180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�J ParagraL     60 ,  0 ,  0 ,  0 , None , !�J Paragraph , Arial ,  10 , M    , None , !�J Paragraph , Arial ,  10 ,  180 ,  250 ,  20 ,N   raph , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0O   ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�J Parag`   20 ,  0 , -1 , -1 , None , !�L Sub Heading , Arial ,  12 , a    60 ,  0 ,  0 ,  0 , None , !�N Mono Spaced , Courier ,  10R   ne , !�N Mono Spaced , Courier ,  10 ,  180 ,  250 ,  20 , S   Courier ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , NoT    250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�N Mono Spaced , U     0 ,  0 , None , !�N Mono Spaced , Courier ,  10 ,  180 , V    Jump Label , Arial ,  10 ,  180 ,  250 ,  20 ,  20 ,  10 ,W     10 ,  180 ,  250 ,  20 ,  20 ,  10 ,  0 ,  0 , None , !�LX    20 ,  20 ,  10 ,  0 ,  0 , None , !�L Jump Label , Arial ,Y   ,  0 , None , !�L Jump Label , Arial ,  10 ,  180 ,  250 , Z   p Label , Arial ,  10 ,  180 ,  250 ,  20 ,  20 ,  10 ,  0 [    ,  180 ,  250 ,  20 ,  20 ,  10 ,  0 ,  0 , None , !�L Jum\    ,  20 ,  0 , -1 , -1 , None , !�L Jump Label , Arial ,  12]    , None , !�L Sub Heading , Arial ,  12 ,  180 ,  250 ,  40^   ding , Arial ,  12 ,  180 ,  250 ,  40 ,  20 ,  0 , -1 , -1_    180 ,  250 ,  40 ,  20 ,  0 , -1 , -1 , None , !�L Sub Heap    ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�N Monoq   10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�R Bib   60 ,  0 ,  0 ,  0 , None , !�Q Bitmap Paragraph , Arial ,  c    !�Q Bitmap Paragraph , Arial ,  10 ,  180 ,  250 ,  20 ,  d   ial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None ,e    20 ,  60 ,  0 ,  0 ,  0 , None , !�Q Bitmap Paragraph , Arf    None , !�Q Bitmap Paragraph , Arial ,  10 ,  180 ,  250 , g   ph , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 ,h    250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�Q Bitmap Paragrai   ,  0 ,  0 ,  0 , None , !�H Footnote , Arial ,  8 ,  180 , j   None , !�H Footnote , Arial ,  8 ,  180 ,  250 ,  20 ,  60 k   te , Arial ,  8 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , l     180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�H Footnom   0 ,  60 ,  0 ,  0 ,  0 , None , !�H Footnote , Arial ,  8 ,n    ,  0 , None , !�H Footnote , Arial ,  8 ,  180 ,  250 ,  2o    Spaced , Courier ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0�   tmap Jump Label , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  �   �R Enumerated Bullet , Arial ,  10 ,  180 ,  250 ,  20 ,  6r   l ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !s    ,  60 ,  0 ,  0 ,  0 , None , !�R Enumerated Bullet , Ariat    ,  0 , None , !�G Bullet , Arial ,  10 ,  180 ,  250 ,  20u   �G Bullet , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0v   l ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !w     250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�G Bullet , Ariax   60 ,  0 ,  0 ,  0 , Box , !�G Bullet , Arial ,  10 ,  180 ,y   0 , None , !�F Bullet , Arial ,  10 ,  180 ,  250 ,  20 ,  z   Label , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  {   ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�R Bitmap Jump |   0 ,  0 , None , !�R Bitmap Jump Label , Arial ,  10 ,  180 }   Jump Label , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  ~    180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�R Bitmap    0 ,  0 ,  0 , None , !�R Bitmap Jump Label , Arial ,  10 , �   0 ,  0 ,  0 ,  0 , None , !�R Enumerated Bullet , Arial ,  �    ,  10 ,  440 ,  250 ,  10 ,  10 ,  0 ,  0 ,  0 , None , !��     10 ,  10 ,  0 ,  0 ,  0 , None , !�M Outline Leaf , Arial�     0 , None , !�M Outline Leaf , Arial ,  10 ,  440 ,  250 ,�   ne Leaf , Arial ,  10 ,  440 ,  250 ,  10 ,  10 ,  0 ,  0 ,�   ,  180 ,  250 ,  10 ,  10 ,  0 ,  0 ,  0 , None , !�M Outli�   0 ,  0 ,  0 ,  0 , None , !�O Outline Branch , Arial ,  10 �   , !�O Outline Branch , Arial ,  10 ,  180 ,  250 ,  10 ,  1�   rial ,  10 ,  180 ,  250 ,  10 ,  10 ,  0 ,  0 ,  0 , None �    ,  10 ,  10 ,  0 ,  0 ,  0 , None , !�O Outline Branch , A�     0 , None , !�O Outline Branch , Arial ,  10 ,  180 ,  250�    Branch , Arial ,  10 ,  180 ,  250 ,  10 ,  10 ,  0 ,  0 ,�    180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�O Outline�   0 ,  0 ,  0 , None , !�R Enumerated Bullet , Arial ,  10 , �   umerated Bullet , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  �   10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�R En�   M Outline Leaf , Arial ,  10 ,  440 ,  250 ,  10 ,  10 ,  0�   tter Label , Arial ,  12 ,  180 ,  250 ,  20 ,  60 ,  0 , -�   180 ,  250 ,  20 ,  60 ,  0 , -1 ,  0 , None , !�S Index Le�   , -1 ,  0 , None , !�S Index Letter Label , Arial ,  12 ,  �    Letter Label , Arial ,  12 ,  180 ,  250 ,  20 ,  60 ,  0 �   ,  180 ,  250 ,  20 ,  60 ,  0 , -1 ,  0 , None , !�S Index�    0 , -1 ,  0 , None , !�S Index Letter Label , Arial ,  12 �   dex Letter Label , Arial ,  12 ,  180 ,  250 ,  20 ,  60 , �   10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�S In�   50 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�E Line , Arial ,  �    ,  0 ,  0 ,  0 , None , !�E Line , Arial ,  10 ,  180 ,  2�   0 , None , !�E Line , Arial ,  10 ,  180 ,  250 ,  20 ,  60�    Line , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  �   ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�E�     250 ,  10 ,  10 ,  0 ,  0 ,  0 , None , !�E Line , Arial �    ,  0 ,  0 , None , !�M Outline Leaf , Arial ,  10 ,  440 ,��   1 ,  0 , None , !�F Index , Arial ,  10 ,  180 ,  250 ,  20�    60 ,  0 ,  0 ,  0 , None , !�I Glossary , Arial ,  10 ,  1�    , None , !�I Glossary , Arial ,  10 ,  180 ,  250 ,  20 , �   abel , Arial ,  12 ,  180 ,  250 ,  20 ,  60 ,  0 , -1 ,  0�   0 ,  20 ,  60 ,  0 , -1 ,  0 , None , !�V Glossary Letter L�   None , !�V Glossary Letter Label , Arial ,  12 ,  180 ,  25�   l , Arial ,  12 ,  180 ,  250 ,  20 ,  60 ,  0 , -1 ,  0 , �     20 ,  60 ,  0 , -1 ,  0 , None , !�V Glossary Letter Labe�   e , !�V Glossary Letter Label , Arial ,  12 ,  180 ,  250 ,�    Arial ,  12 ,  180 ,  250 ,  20 ,  60 ,  0 , -1 ,  0 , Non�   0 ,  60 ,  0 ,  0 ,  0 , None , !�V Glossary Letter Label ,�    0 ,  0 , None , !�F Index , Arial ,  10 ,  180 ,  250 ,  2�   , !�F Index , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 , �   rial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None �   80 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�F Index , A�    ,  60 ,  0 ,  0 ,  0 , None , !�F Index , Arial ,  10 ,  1�   80 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�I Glossary �   ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�D Bar ,�    ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�D Bar , Arial ,  10 �   ,  0 ,  0 ,  0 , None , !�D Bar , Arial ,  10 ,  180 ,  250�   0 , None , !�D Bar , Arial ,  10 ,  180 ,  250 ,  20 ,  60 �   D Bar , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  �    ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !��     250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�F Image , Arial�   60 ,  0 ,  0 ,  0 , None , !�F Image , Arial ,  10 ,  180 ,�    0 , None , !�F Image , Arial ,  10 ,  180 ,  250 ,  20 ,  �    Image , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 , �   ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�F�    250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�F Image , Arial �     0 ,  0 ,  0 , None , !�I Glossary , Arial ,  10 ,  180 , �   ne , !�I Glossary , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,�   , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , Noj�    Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , Non�   ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,�   1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  �   e , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !��   !�;  , Arial ,  10 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 , Non�    ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , �   0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0�    0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  �   ,  0 ,  0 ,  0 , None , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 , �    ,  0 ,  0 , None , !�;  , Arial ,  10 ,  0 ,  0 ,  0 ,  0 �   ne , !�F Table , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0�   , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , No�     180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�F Table �    20 ,  60 ,  0 ,  0 ,  0 , None , !�F Table , Arial ,  10 ,�   ,  0 ,  0 , None , !�F Table , Arial ,  10 ,  180 ,  250 , �   e , !�F Table , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 "�     0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�;  , Arial ,  10 ,�    0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 , None , !�1  ,  ,  0 ,  0�    0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�;  , Arial ,  10 , �     0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 , �     ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,�    , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1�   �;  , Arial ,  10 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 , None�   ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�    ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 �   0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0�     0 ,  0 ,  0 , None , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  �     0 ,  0 ,  0 ,  , !�;  , Arial ,  10 ,  0 ,  0 ,  0 ,  0 ,�   ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,�    ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 �   0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0�     0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 , None , !�1  ,  ,  0 ,  ��    ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 �   e of the INIVISICLUES was to provide hints to several parts�   ch the idea of interactive providing hints. The main purpos�   ersions of the INVISICLUES(TM), but plane text does not mat�   inally the purpose of this software was to renew the INVISI�   CLUES(TM) in an electronical way to prevent the final loss �   of information. In addition there are different places in t�   he internet where you can find more or less complete text vm  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�   y /Popup /Just L /Text !�C /L /Jump Referenzen /Link /Macro�    THL software and THL files ?!�1 /L /Jump /Link /Macro /Pla�   192,192), 0!�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  9   	  � 1000   �  ��7j     � Contents;Overview;�� B�       0 ,  0 ,  0 ,  , !�                                       �     0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 , �   ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,    of a game. These hints were divided into different topics   or further information.����Please remember: The sole intent�   vide additional language support packs. Please contact me f�    help. I would be very pleased if anyone out there will pro�   ble shall be supported by the user interface and the online�   avaible to a wide range of users as many languages as possi�   . (This is not limited to games !).��To make this software �   is project and develop their favourite hints to other users�   file collection. And everyone is invited to take part in th�    the new purpose of The Hint Library is to build up a hint �   lso the capabilities to create new hint collections. By now�   stem I decided not just to provide a read-only system but a�   elp as you need or as you wish. ����While developing the sy�   on with text-based solutions is that you just get as much h�   vided. The main advantage of these collections in comparisi�   while the hints were sorted due to the level of details pro�   of this software is collecting information, It must not be  ur raw data is invisible. ��Information about compiling you  ion.��The compiler part, which generates a THL file from yo  n on creating THL files please refer to The THL Editor sect  P, JPEG, TARGA, PCX) in your files.��For further informatio  text, multimedia files ( Sound, Videos ), and pictures ( BM  collections with an easy to use interface. You can include   editor, which provides capabilites for creating new hint   e refer to Read THL-Files section.��The second part is the 	  a files( e.g. MIDI, AVI,...)��For further information pleas
  he following types of hints: Text, pictures, and  multimedi  receiving  of information shall be avoided. You will meet t   know explicitly requested information only. Inadvertandly   , provides capabilites for browsing hintfiles. You will get  Mainly there are two sections. The first one, ther Reader   used for any commercial purposes.����About the software:��    can find in Creating own THL files section.����Please send!  lay  PCX-,TGA- and JPEG-Files. Contact:��Meister@rz.fhtw-be  ef Meister. Partially his MPICVIEW-Project is used to disp  :����Beta-Testers:��Klaus Meier��Alen Tomasic����Detl  �  	  � 2000   �  ��;�   :  �5 Hint files;Infocom;Lang  uage files;Languages;Overview;�� F�     � Introduction  �� U�     �  �� 	��  �
-�   !�* /T /Just L /Text Intro�   duction and Overview!�
 /N /Just L!��
/P /Just L /Text Orig  �    �    �  ��;�   1  �, Author;Borland Delphi;Greet  ings;Information;�� B�     � Credits�� Q�     �  ��   	�}  �-�   !� /T /Just L /Text Credits!�
 /N /Just L!�  �/P /Just L /Text Author: Stefan Meier����Special thanks �  ag /Link /Macro /Play /popup /Just L /Text License Agreemen   /Play /popup /Just L /Text Credits!�P /L /Jump Lizenzvertrw  n Meier, Erfstr. 65, 52249 Eschweiler��AOL:      SMeier7777   questions, announces or bug reports to:��Mail:       Stefaj0  rlin.de����All former Infocom programmers, which made their#   of the notice.  Termination of the right to distribute doe$  s not affect distributors' other duties in this license.���%  �Many thanks go to Detlef Meister for his freeware project &  MPICVIEW. Parts of this project are used for displaying JPE'  G,TARGA and PCX files.��You can contact Detlef Meister at:�(  �Meister@rz.fhtw-berlin.de�� ��Enjoy The Hint Library!����C)  ontact:��Stefan Meier, Erfstr. 65, D-52249 Eschweiler, Germ*  any��AOL:��SMeier7777��E-Mail:��SMeier7777@aol.com��Stefan.    Meier@post.rwth-aachen.de��  
� �                        �    ���� 
V 0 7 P     � Topic@Lizenzvertrag  �    �  �H�� 
 - 4 M     � Topic@Einleitung  �      �  4��� 
 - 4 I     � Topic@Referenzen  �                                                                   .  Library 1.0 was created using Borland Delphi 2.0.��  
� �/   adventures a milestone in computer history.������The Hint ""   must stop distributing this archive 30 days after the date3  e to the ftp-Site given at the bottom of this document.����4  Distribution through retail and wholesale stores requires s5  pecific written permission.��Distribution through "magazine6  - compact disks" or "magazines-floppy disks" requires speci7  fic written permission.��No distributor may charge more tha8  n $8 US (or the appropriate value in other currencies, e.g.9   12 DM) for this archive.����Vendors' entire collection of :  THL files must be stored on a reasonably small number of di;  sks; distribution of hint files over excessive numbers of d<  isks is prohibited.  No more than $8 US (or the appropriate=   value in other currencies, e.g. 12 DM) may be charged for >  any disk containing THL files.��These terms are a condition?   of distribution of this archive and apply to all THL files@   written by any hint author.����Right to distribute this ar1  chive may be terminated by written notice, and distributors�2  ase send a copy to me. The easiest way is to upload the filC   documentation are provided "AS IS" and without warranty ofD   any kind and the author expressly disclaims all other warrE  anties,��express or implied, including, but not limited to,F   the implied warranties of merchantability and fitness for G  a particular purpose. Under no circumstances shall Stefan MH  eier be liable for any incidental, special or consequentialI   damages that result from the use or inability to use the sJ  oftware or related documentation, even if Stefan Meier has K  been advised of the possibility of such damages.����If you L  intent to write THL-files with the included editor and distM  ribute them you should always contact me to tell me about yN  our project and check out if anyone else is working on a hiO  nt file for the given game. Although the use of the softwarP  e is free you are NOT ALLOWED to take charge for your indivA  idual THL-files.  If you want to spread your THL-Files, ple�B  is software in your possession.����The software and relatedS  ement between you and Stefan Meier covering your use of TheT   Hint Library. Be sure to read the following agreement befoU  re using the software. IF YOU DO NOT AGREE TO THE TERMS OF V  THIS AGREEMENT, DO NOT USE THE SOFTWARE AND DESTROY ALL COPW  IES OF IT.��This copyright software is distributed as freewX  are. You may use this software without any charge and may dY  istribute to others. The software is owned by Stefan Meier Z  and is protected by FR Germany copyright laws and internati[  onal treaty provisions. Therefore, you must treat the softw\  are like any other copyrighted material (e.g., a book or mu]  sical recording).����You may not rent or lease the software^  , nor may you modify, adapt, translate, reverse engineer, d_  ecompile, or disassemble the software.��If you violate any `  part of this agreement, your right to use this software terQ  minates automatically and you then destroy all copies of thR  ment!�
 /N /Just L!�(/P /Just L /Text This is a legal agreq  ing your own files.!�h /R /Link E:\WORK\HINT_R~1\HELPFILE\Eb  tion of THL files you can find at: The THL editor and Creatc  a new file. Information on editor instructions and the cread  NEWFILE.BMP /Just L /Text Open the THL editor for creating e  es of the THL files.!�� /R /Link E:\WORK\HINT_R~1\HELPFILE\f  n verbose mode. You will not see the filenames but the titlg  HINT_R~1\HELPFILE\VOPEN.BMP /Just L /Text Open a THL file ih  ou cam find in the THL Reader section.!�� /R /Link E:\WORK\i   THL file for reading hints. Information on reading hints yj   E:\WORK\HINT_R~1\HELPFILE\OPENBTN.BMP /Just L /Text Open a�  �  ���� 
m - 4 I     � Topic@Referenzen  �    �   !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�o    �  	  � 7000   �  ��>�   +  �& Conditions;License;Dp  istribution rules;�� I�     � Licence Ageement�� X�  a     �  �� 	�&  f-�   !�" /T /Just L /Text License Agree��  XISTF~1.BMP /Just L /Text Open an existing THR file with th�  ing the file to edit.��!��/R /Link E:\WORK\HINT_R~1\HELPFIr  e opens the editor and brings up a file open box for chooss  editor window with a blank formular��Editor - Edit hintfilt  BMP /Just L /Text Editor - Create new hintfile opens the u  ibrary��!�� /R /Link E:\WORK\HINT_R~1\HELPFILE.GB\EDITOR~1.v  by title and opening the Reader..��Exit exists The Hint Lw  the Reader.��Select Verbose open for choosing a THL file x  ext Select File open for choosing a THL file and opening y   /Link E:\WORK\HINT_R~1\HELPFILE.GB\DATEIM~1.BMP /Just L /Tz  int Library!�& /H 2 /Just L /Text The program menues:!�� /R{  E:\WORK\HINT_R~1\HELPFILE\EXIT.BMP /Just L /Text Exit The H|   like program version and contact information.!�O /R /Link }  ~1\HELPFILE\INFO.BMP /Just L /Text Show program information~  ust L /Text Open this help file.!�� /R /Link E:\WORK\HINT_R  e editor.!�N /R /Link E:\WORK\HINT_R~1\HELPFILE\HELP.BMP /J"�  LE.GB\SPRACH~1.BMP /Just L /Text Use Language - Select lan�  ��/R /Link E:\WORK\HINT_R~1\HELPFILE.GB\HILFEM~1.BMP /Just�    	  � 3000   �  ��:x   "  � Main window;Menues;Langu�  ages;�� E�     � Operating instructions�� T�     �  �  �� 	��
  C
-�   !�' /T /Just L /Text Operating instructio�  ns!�
 /N /Just L!�Y /P /Just L /Text After starting The Hin�  t Library you will encounter the following window:!�6 /I /L�  ink E:\WORK\HINT_R~1\HELPFILE.GB\MAIN.BMP /Just L!� /H /Juk  st L /Text !�  /H 2 /Just L /Text Speedbuttons:!�� /R /Link�  nguage will be selected each time you start automatically.!�  ge - Save language setting you can decide if the chosen la�  language packages please refer to THL homepage. WithLangua�  ded, but the system can easily be extended. For additional �  kage. By default only the English language package is inclu�   �  �.�� 
� ) 0 I     � Topic@Inhalt  �    �  �  guage to open a dialog for choosing a language support pac"�   L /Text Use Help - Contents to start online help and go �     !� /T /Just L /Text THL-Dateien!�
 /N /Just L!�/P /J�  �     � What�s a THL-File ?�� ^�     �  �� 	�G  a-��  eien;Hinweise;Bilder;Formate;THL-Dateien;THR-Dateien;�� O�  ..  �    �    �    �  ��H�   H  �C Multimedia-Dat�  L!�r /L /Jump Was sind THL Dateien... /Link /Macro /Play /p�    �-�   !� /T /Just L /Text The THL editor!�
 /N /Just �  iles,edit;�� F�     �
 The editor�� U�     �  �� 	�G�  �  	  � 5000   �  ��;}   &  �! Editor;THL Editor;THL f�    	  � 3000   �  ��:x   "  � Main window;Menues;Langu                                                                   act adresses and other usefull information.  
� �        �  rmation dialog where you can find the program version, cont�   on using the Windows help system��Info brings up an info�  es by key words��Help - Using help shows you instructions�  to contents page��Use Help - Search to search the helpfil�  T  ���� 
� : A V   "  � Topic@Was sind THL Dateien.�  ace.!�9 /B /Just L /Text Compile the editor data into a THL�  r anymore. Always keep a copy of your THR-File at a save pl�  .��CAUTION: THL-File can not be edited with the THL-Edito�  ommened). A THR-File saves your data without compiling them�  t L /Text Eventually save your data as THR-File (highly rec�  hints, include pictures, ... with the THL-Editor!�� /B /Jus�  es consists of three main steps:!�G /B /Just L /Text Enter �  or ordinary texteditors. In general the creation of THL-Fil�   the "reader" of this software, but they are not suitable f�  ures and multimediadata. They are designed for the use with�  L /Text THL-Files are binary files which contain text, pict�   !� /T /Just L /Text THL-Files!�
 /N /Just L!�/P /Just �      � What�s a THL-File ?�� ^�     �  �� 	�K  g-�  �  formats;Hints;Multimedia files;THL files;THR files;�� O� �  ..  �    �    �    �  ��H�   F  �A Pictures;File ��  -File.!� /H 1 /Just L /Text !�2 /H 1 /Just L /Text The str�  opup /Just L /Text What are THL files, how are they created�  s 1..6����Invalid structure:��Topic1 ---> Hints 1..3��Topic�  Topic2 ---> Subtopic1, Subtopic2��Topic3 ---> Picture, Hint�  t Two examples:��Valid structure:��Topic1 ---> Hints 1..3���  t recommened due to compability reasons.!�� /P /Just L /Tex�  V. Some additional formats are supported, but the use is no�  Text Multimedia-Files, suported formats: WAV, AVI, MIDI, MO�  ctures and attach independent descriptions.!�� /B /Just L /�  g, PCX, Targa��Special features: You may define parts of pi�  /Just L /Text Pictures, supported file formats: Bitmap, JPe�  2 /B /Just L /Text Text ( single or multiple lines )!�� /B �  e combined at one level.��There are different hint types:!��  ther contain subtopics or hints. Hints and topics can not b�  t collection is divided into deveral topics. These topic ei�  ucture of THR/THL-Files:!�� /P /Just L /Text Ordinary a hin�  ?!�u /L /Jump Eigenentwicklung von Hinweissammlungen /Link �  any copyrights. Ordinarily it is prohibited to transform co�  mmercial hint books into electronical systems. If you have �  doubt about legimitation please contact the author of the o�  riginal.!�� /B /Just L /Text You should spread THL files on�  ly. Remember that anyone is able to edit the data in a THR �  file, but always keep a copy of your THR file at a secure p�  lace. A THL file can not be edited with the THL editor.!��  /B /Just L /Text Please send a copy of your THL file to me.�  ng ftp-site:��ftp://members.aol.com/thlhome/incoming��Alt�  ernativly you can send the file by mail or name a internet     site where I can download the file.  
� �                �   The easiest way to do is uploading the file to the followi�  P  �W�� 

 - 4 M     � Topic@Der Editor  �    4  les.!�k /L /Jump Die Bedienung des Editors /Link /Macro /Pl�  /Macro /Play /popup /Just L /Text Development of own THL fij�  sions.!�� /B /Just L /Text Please make sure not to violate �  Hinweissammlungen  �    �    �    �  ��W�   -  �(�   Userdefined files;Development;THL files;�� ^�   !  � Cr�  eation of hint collections�� m�     �  �� 	��  �-�  	�   !�, /T /Just L /Text Creating your own THL files!�
 /N /Ju�  st L!�v /P /Just L /Text If you wish to design and spread o�  wn hint collections, please pay attention to the following �  advices:!� /B /Just L /Text Before starting your work you �  should contact me to check if anyone else is working on a f�  ile about your topic. This is done to avoid double works on�   one topic and to make it possible to me to keep an eye on �  the progress of the THL project.!�� /B /Just L /Text Think �  about the structure of your hint collection. Where can ques�  tions occur ? When is picture support usefull ? Which logic�  al parts can be defined ?!�_ /B /Just L /Text Compare your �  solution with different solutions to prevent errors or omis��  �  �^�� 
 I P e   1  �, Topic@Eigenentwicklung von �  /Text Where can I get... ?!�
 /N /Just L!�� /B /Just L /Tex�   I get...?�� X�     �  �� 	��  � -�   !�% /T /Just L �  ks;New program versions;THL files;�� I�     � Where can�    �  	  � 8000   �  ��>�   ;  �6 Language support pac�  �  ��� 
 0 7 P     � Topic@Wo gibt es...  �  �  �  �E�� 
� 0 7 P     � Topic@Wo gibt es...  �  `    !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  t!�; /P /Just L /Text ������The Hint Library � 1996 Stefan �    �  	  � 7000   �  ��>�   8  �3 Benutzung, Bedingung�  [  V�� 
| 0 7 P     � Topic@Lizenzvertrag  �  n  /  #��� 
 0 7 P     � Topic@Lizenzvertrag  �  �   Entwicklung;Eigene Dateien;THL-Dateien;�� ^�   +  � Cre�  ation of hint collectionsammlungen�� m�     �  �� 	���    �-�  	 !�0 /T /Just L /Text Entwicklung eigener THL-Date�  ien!�
 /N /Just L!�� /P /Just L /Text Wenn Sie beabsichtige"�  t New program versions, language support packages, and THL �  xt This button opens a Save File-Dialog for saving your pro�  ject as THR file. You need this THR file for later changes.�   It is highly recommend to save THR files of each important�   development state of your project.!�C /E /Just L /Text Thi�  s button compiles your project into a THL file.!�j /E /Just�  P  V��� 
s : A V   "  � Topic@Was sind THL Dateien.�  Hinweissammlungen  �    �    �    �  ��W�   ,  �'�   L /Text Press this button to exit THL Editor. Always save     your project before leaving the editor.  
           ?  N  ΍�� 
� < C \   $  � Topic@Die Bedienung des Edi�    ^��� 
	 , 3 L     � Topic@Bedienung  �    �k    	  � 3000   �  ��:w   �� � Main window;Menues;Langu�  Z  5��� 
� , 3 L     � Topic@Bedienung  �    �    Meier  
� �                                                   !�                                                        "�  dditional information about your project.!�� /E /Just L /Te  n delete all children of this entry. Use this function care  fully !!�� /E /Just L /Text This buttons moves the currentl  y selected item within its level upwards. Associated childr  en will be moved either.!�$ /E /Just L /Text Moving downwar  ds...!�� /E /Just L /Text Enter a title for your document h  ere. This is not a file name, but a title which appears as 	  header in the Reader. This entry is nessesary for successfu
  ll compilation.!�/E /Just L /Text With this button you ca  n choose a font which will be used with the Reader to displ  ay the title of your document. Please note that the use non   standard fonts may cause unwanted  effects on computer sys  tem which do not have the fonts installed.!�� /E /Just L /T  ext Use this window to enter copyright notice, e.g. Writte  n 1996 by Harry Hummel. This field must be filled in for p  roper compilation.!�N /E /Just L /Text Here you can enter a  lete the currently selected entry. Please note that you eve  ecome enabled or disabled.!�[ /E /Just L /Text Pressing thi  s button open a window for adding a new topic to your proje  ct.!�= /E /Just L /Text Here you can add a new hint to your   project.!�� /E /Just L /Text This button opens the picture   editor which is used to add new picture links or area defi  nitions to your project.!��/E /Just L /Text Pressing butto  n no 5 open a window for adding multimedia files to your pr  oject. Please note that normally video files are rather lar  ge and therefore the size of the THL file will increase sig  nificantly. Although the multimedia support of THE HINT LIB  RARY only depends on the capabilites of your system, unusua  l files formats may not be supported by different systems.!  �� /E /Just L /Text Edit the selected entry. The software w   ill select the appropriate window for the entry. It is not   possible to change type of an entry.!�� /E /Just L /Text De�  try. According to your avaible selections the buttons 2-5 b#  tors  �    �  	  � 6000   �  ��J�   |  �w Author;P$  ictures;Edit files;Editor;File formats;Hints;Multimedia fil%  es;Font;Topics;THL files;THL Editor;THR files;Title;�� U&      � Using the THL editor�� d    �  �� 	��  �-�'     !�% /T /Just L /Text Using the THL editor!�
 /N /Just L(  !�R /I /Jump /Link E:\WORK\HINT_R~1\HELPFILE.GB\EDITOR.BMP )  /Macro /Play /Popup /Just L!�L /P /Just L /Text PLEASE PAY *  ATTENTION TO THE ADVICES ON CREATING THL FILES !!��/E /Jus+  t L /Text This tree view shows your current project. Hints ,  are marked with the prefix HINT, pictures are marked with P-  IC, and multimedia files are marked with MM. You always wil.  l see the starting characters of a title. The root director/  y contains topics only. Topics either contain subtopics or 0  hints, pictures, or multimedia files. When adding new entri!  es the currently selected entry becomes owner of the new en�"  �  M��� 
 < C \   $  � Topic@Die Bedienung des Edi3  f you close this window with the OK button, the new topic w    ill be added to your project.  
� �                      �  ay /popup /Just L /Text Instructions on using the editor  z  , Bedienung;Editor;�� U%    � Using the THL editortor5  s�� d5    �  �� 	�  |-�   !�% /T /Just L /Text Usi6  ng the THL editor!�
 /N /Just L!�O /I /Jump /Link E:\WORK\H7  INT_R~1\HELPFILE\EDITOR.BMP /Macro /Play /Popup /Just L!�P 8  /P /Just L /Text BITTE BEACHTEN SIE DIE HINWEISE ZUM ERSTEL9  LEN VON THL-DATEIEN !!�^/E /Just L /Text Hier sehen Sie Ih:  r Projekt als Baumansicht, Hinweise enthalten vor ihrem Ein;  trag das Schl�sselwort HINT, Bilder das Schl�sselwort PIC u<  nd Multimediadateien MM. Bei Themen sehen Sie sie ersten Bu=  chstaben des Titels. Das Hauptverzeichnis (<<<Script>>>) ka>  nn nur Themen enthalten. Die einzelnen Themen enthalten ENT�  �  y
�� 
� 9 @ Y   !  � Topic@Das Multimedia Fenste2  t L /Text Enter the title of your topic at the TEXT line. IC  nster  �    �  	  � 5020   �  ��K�     � Hint;AdD  ding hints;Text;�� V�     � The hint edit window�� e�E       �  �� 	��  %-�   !�% /T /Just L /Text The hint edF  it window!�
 /N /Just L!�T /I /Jump /Link E:\WORK\HINT_R~1\G  HELPFILE.GB\HINTEDIT.BMP /Macro /Play /Popup /Just L!�� /P H  /Just L /Text Enter your text into the Text field. If you cI  lose the window with the OK button the new hint will be add    ed to your project.  
� �                                K  �  X��� 
� < C \   $  � Topic@Das Themen EditierfenL  ster  �    �  	  � 5030   �  ��J~     � Text;AddM  ing topics;�� U�     � The topic edit window�� d�   N    �  �� 	��  3-�   !�& /T /Just L /Text The topic edit P  window!�
 /N /Just L!�S /I /Jump /Link E:\WORK\HINT_R~1\HEL_  r>!�1 Bild-Editierfenster,Das Bilder Editierfenster, 0,!�S A  PFILE.GB\TOPEDIT.BMP /Macro /Play /Popup /Just L!�� /P /Jus�  ,(Global), 0,<Das Multimedia Fenster>!�+ Read THL-Files,(Gla  escription. On selecting a new picture the complete pictureR  e added to the hotspot list. Now you just have to enter a dS  . On releasing the left mouse button the marked area will bT   into the picture and marked the area by dragging the mouseU  eparate picture areas: Click and hold the left mouse buttonV  ename at the FILE field. Use the hotspot editor to define sW  /Play /Popup /Just L!��/P /Just L /Text Please enter a filX  Jump /Link E:\WORK\HINT_R~1\HELPFILE.GB\PICEDIT.BMP /Macro Y  /Just L /Text The picture edit window!�
 /N /Just L!�S /I /Z  icture edit window�� d�     �  �� 	�A  f-�   !�( /T [  ordinates;Pictures;Progress indicator;�� U�     � The p\  ster  �    �  	  � 5010   �  ��J�   3  �. Areas;Co]  J  c�� 
� < C \   $  � Topic@Das Bilder Editierfenh  Creating own THL files section,(Global), 0,<Eigenentwicklun�  �  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  p   will be added to the hotspot list automatically. Show shouc   L /Text The multimedia edit window!�
 /N /Just L!�R /I /Jud  mp /Link E:\WORK\HINT_R~1\HELPFILE.GB\MMEDIT.BMP /Macro /Ple  ay /Popup /Just L!�� /P /Just L /Text Please enter a filenaf  me in the File field or choose a file with the Browse buttog  n. Afterwards enter a description f�r the multimedia hint a�  t the descriptiion field. Closing the window with the OK bu}  g von Hinweissammlungen>!� CREATING THL FILES,(Global), 0,�  ster  �    �  	  � 5010   �  ��J�   3  �. Areas;Pii  ctures;Progress indicator;Coordinates;�� U�     � The pj  �  x�� 
� , 3 L     � Topic@Bedienung  �    �    rate entries for the THL files.  
� �                    l  er picture in your project, the compiler will generate sepam  o your project. Although you only will see a single entry pn  he window with the OK button, the new entry will be added to  ld edit the description or remove the item.��If you close t"b  a edit window�� h�     �  �� 	�r  �-�   !�+ /T /Just�  Hinweisdateien;Infocom;�berblick;�� F�     � Introductir  on�� U�     �  �� 	��  �-�   !�* /T /Just L /Text In    thlhome/index.htm����Enjoy THE HINT LIBRARY !��  
� �    t  tp://members.aol.com/thlhome��oder��http://members.aol.com/u  .Meier@post.rwth-aachen.de����The Hint Library Homepage:��fv  ��e-Mail:   SMeier7777@aol.com oder��                Stefan�  nweissammlungen>!�N ERSTELLEN VON THL-DATEIEN,(Global), 0,<x   THL-Dateien erstellen,(Global), 0,<Eigenentwicklung von Hi�  rmate;Dateien bearbeiten;THL-Dateien;THR-Dateien;THL-Editory  ditor>!�' Der-THL-Editor,(Global), 0,<Der Editor>!�Q Eigene{  von Hinweissammlungen>!�' Der THL-Editor,(Global), 0,<Der E|  !�M Creating your own files.,(Global), 0,<Eigenentwicklung   {  ���� 
� @ G `   (  �# Topic@Das Multimedia Editie�  rfenster  �    �  	  � 5040   �  ��N�   '  �" Fileq   description;Multimedia files;�� Y�     � The multimedi��  �  	  � 2000   �  ��;�   =  �8 Sprachdateien;Sprachen;�  Jump /Link E:\WORK\HINT_R~1\HELPFILE.GB\READER.BMP /Macro /�  Play /Popup /Just L!�� /P /Just L /Text The list box centre�  d in the window displays the main topics contained in the f�  ile. Double-clicking an item opens the specific topic. Ther�  e will will either encounter different subtopics or hints:!�  �� /R /Link E:\WORK\HINT_R~1\HELPFILE.GB\HINTPIC.BMP /Just �  L /Text Text hints: Double-clicking a hint item opens the h�  int window. Because hints are sorted to their level of deta�  il a warning will raise if you try to read hint no 3 before�   hint no 2.!�� /R /Link E:\WORK\HINT_R~1\HELPFILE.GB\MMPIC.�  BMP /Just L /Text Multimedia hints: Double-clicking a multi�  media item brings up a multimedia control panel..!�� /R /Li�  nk E:\WORK\HINT_R~1\HELPFILE\PICPIC.BMP /Just L /Text Pictu�  re hints: Double-clicking a picture item opens the picture     display window.  
� �                                    ��  a THL file you will encounter the following window:!�R /I /�  edia files;Multimedia contral;Multimedia player;�� R�   !�  r  �    �  	  � 4030   �  ��G�   @  �; Play multim�  Eigenentwicklung von Hinweissammlungen>!�8 Hinweis-Anzeigef�  ende Fenster. If you decide not to read the hiont yet, you �  can abort by pressing the Close icon in the upper right cor    ner.  
� �                                               �  =  ��� 
� 6 = V     � Topic@Das Hinweis Fenster�    �  	  � 4000   �  ��?�   &  �! Hinweise lesen;THL-    bers.aol.com/thlhome  
� �                                   !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�             �  �  ��� 
 1 8 Q     � Topic@Der THL Reader  �  �    �  	  � 4000   �  ��?}   "  � Read hints;Reader;T�  HL Reader;�� J�     � The THL Reader�� Y�     �  ���   	��  �-�   !� /T /Just L /Text The THL Reader!�
 /N /J�  ust L!�e /P /Just L /Text After opening and compilation of ��    � The multimedia control panel�� a�     �  �� 	�.  �  EW.BMP /Macro /Play /Popup /Just L!��/P /Just L /Text Afte�  r selecting a hint you will encounter the following window.�   For reading the hint you have to click the SHOW HINT butto�  n. After reading the hint you can close the window by presi�  ng the close button. This hint will be marked as "read". ���  Wenn Sie einen Hinweis ausgew�hlt haben, sehen Sie das folg�  -lesen,(Global), 0,<(None)>!�5 Hinweis-Editierfenster,Das H�  enster,(Global), 0,<Das Hinweis Fenster>!�* Hinweis-Dateien@  r  �    �  	  � 4030   �  ��G�   G  �B Multimedia-    stops a currently running media  
� �                    �  nel is shown. Pressing the OK button closes the window and �   After selecting a multimedia hint the following control pa�  \MMVIEW.BMP /Macro /Play /Popup /Just L!�� /P /Just L /Text�  
 /N /Just L!�R /I /Jump /Link E:\WORK\HINT_R~1\HELPFILE.GB�  D-�   !�- /T /Just L /Text The multimedia control panel!��  ust L!�T /I /Jump /Link E:\WORK\HINT_R~1\HELPFILE.GB\HINTVIB  �  �N�� 
� = D ]   %  �  Topic@Das Hinweis Editierfe�  (  e�� 
� < C \   $  � Topic@Das Bilder Editierfen�    D��� 
� : A Z   "  � Topic@Das Bildanzeige Fenst�  er  �    �  	  � 4010   �  ��H�   !  � Pictures;P�  rogress indicator;�� S�     � The picture display windo�  w�� b�     �  �� 	�  =-�   !�+ /T /Just L /Text The�   picture display window!�
 /N /Just L!�S /I /Jump /Link E:\�  inweis Editierfenster, 0,!�; Multimedia-Editierfenster,Das �  WORK\HINT_R~1\HELPFILE.GB\PICVIEW.BMP /Macro /Play /Popup /�  Just L!�� /P /Just L /Text The progress indicator in the lo�  wer left corner shows refers to the file loading process. P�  ressing the Close button exists the display window.  
� ��    �    �  	  � 4020   �  ��D{     � Hidden hint;Sh�  ow hint;�� O�     � The hint window�� ^�     �  �� �  	��  J-�   !�  /T /Just L /Text The hint window!�
 /N /J�    ���� 
� 6 = V     � Topic@Das Hinweis Fenster�  (Global), 0,<Der THL Reader>!�- THL-Homepage nach,(Global),�  Editierfenster,Das Themen Editierfenster, 0,!�' THL Reader,�  ader>!�' The THL editor,(Global), 0,<Der Editor>!�3 Themen-�  obal), 0,<Der THL Reader>!�# Reader,(Global), 0,<Der THL Re+  �  [��� 
n 0 7 P     � Topic@Wo gibt es...  �      2 ---> Subtopic1, Hints1..9 ( ERROR )��...  
� �         l  �  ���� 
l 0 7 P     � Topic@Lizenzvertrag  �  s  �  ���� 
� I P e   1  �, Topic@Eigenentwicklung von �  �  ���� 
� < C \   $  � Topic@Die Bedienung des Edi�  tors  �    �  	  � 6000   �  ��J�   �  �� Schrifta�  rt;Autor;Titel;Themen;Bilder;Multimedia-Dateien;Hinweise;Fo�  �  <��� 
� 1 8 Q     � Topic@Der THL Reader  �      
� �                                                      �  7  ���� 
� 9 @ Y   !  � Topic@Das Multimedia Fenste    tton adds the new entry to your project.  
� �                0,<Wo gibt es...>!�                                                                                                      �                                                             �  files:��http://members.aol.com/thlhome/index.htm��ftp://memQ  Multimedia Editierfenster, 0,!�? Multimedia-Kontrollfenster�  T  ķ�� 
� - 4 M     � Topic@Einleitung  �    �  �  	  � 2000   �  ��;�   =  �8 Sprachdateien;Sprachen;�  Hinweisdateien;Infocom;�berblick;�� F�   �� � IntroduL �   �� U�     �  �� 	�C  z-�   !�) /T /Just L /Text Einl�  eitung und �berblick!�
 /N /Just L!�5/P /Just L /Text Ursp�  r�nglich war dieses Programm nur dazu gedacht, die INVISICL�  UES(TM) zu den alten INFOCOM-Adventures in elektronischer F�  orm wiederaufzubereiten, um zu verhindern, da� diese Inform�  �  ^M�� 
� - 4 M     � Topic@Einleitung  �    �  �  �� 
d , 3 L     � Topic@Bedienung  �    ��  �  nn�� 
� , 3 L     � Topic@Bedienung  �    �